`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:30:16 01/05/2017 
// Design Name: 
// Module Name:    Final 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Final(
	input rst,
	input clk,
	input PSCLK,
	input PSDATA,
	output R,
	output G,
	output B,
	output hsync,
	output vsync
    );

//////////////////////////////////////////////////////////////////////////////////
// Parameter
//////////////////////////////////////////////////////////////////////////////////
//parameter PERIOD = 3000000;

parameter leftX   = 104;
parameter rightX  = 904;
parameter centerX = 504;
parameter topY    = 20;
parameter downY   = 632;

parameter wallW = 20;
parameter hp = 80;
parameter radius = 20;
parameter bInitX = 700;
parameter bInitY = 400;
parameter bStepX = 10;
parameter bStepY = 10;
//parameter StepXinit = 10;
//parameter StepYinit = 10;
//parameter MaxSpeedX = 50;
//parameter MaxSpeedY = 50;
//parameter barAx = 140;
//parameter barBx = 850;
//parameter barL = 100;
parameter barW = 20;
parameter MAX = 10000;

parameter poX = 300;
parameter poY = 200;

// bar
parameter initAX = 140;
parameter initBX = 850;
parameter initY = 300;
parameter uStepX = 20;
parameter uStepY = 20;
parameter leftAX = 140;
parameter rightBX = 850;

//////////////////////////////////////////////////////////////////////////////////
// Wire or Reg
//////////////////////////////////////////////////////////////////////////////////
reg [20:0] x, y;
wire [10:0] vis;
reg nState, cState;
reg [21:0] kReg;
reg [7:0] kData;
reg [3:0] kCounter;
wire check;
reg [30:0] counter;
//reg [4:0] time2;
reg timer;
reg isStop;

// keyboard
reg sig_f0;
reg up, down, right, left, w, s, a, d, sp;

reg [20:0] barAx, barBx;

// speed
//reg [20:0] bStepX, bStepY;
reg [30:0] PERIOD;
//reg [30:0] ppp;

// color
wire black, white;
reg mod1, mod2, mod3;

// object
reg barA, barB;
reg ball;
reg topWall, downWall, leftWall, rightWall;
wire wall;
reg [6:0] barL;
reg cLine;

// Center
reg [10:0] bCenterX, bCenterY;
wire [10:0] pCenterX, pCenterY;
reg bXd, bYd;

// keyboard
reg [30:0] barAy, barBy;

// final
reg aW, bW;
reg Awins, Bwins;
wire [400:0]  B0, B1, B2, B3, B4, B5, B6, B7, B8, B9, B10, B11, B12, B13, B14, B15, B16, B17, B18, B19, B20, B21, B22, B23, B24, B25, B26, B27, B28, B29, B30, B31, B32, B33, B34, B35, B36, B37, B38, B39, B40, B41, B42, B43, B44, B45, B46, B47, B48, B49, B50, B51, B52, B53, B54, B55, B56, B57, B58, B59, B60, B61, B62, B63, B64;
wire [400:0]  A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14, A15, A16, A17, A18, A19, A20, A21, A22, A23, A24, A25, A26, A27, A28, A29, A30, A31, A32, A33, A34, A35, A36, A37, A38, A39, A40, A41, A42, A43, A44, A45, A46, A47, A48, A49, A50, A51, A52, A53, A54, A55, A56, A57, A58, A59, A60, A61, A62, A63, A64, A65, A66, A67;

//////////////////////////////////////////////////////////////////////////////////
// C C
//////////////////////////////////////////////////////////////////////////////////
assign hsync = ~( (x >= 919) && (x < 1039) );
assign vsync = ~( (y >= 659) && (y < 665) );
assign vis = ( (x >= 104) && (x < 904) && (y >= 23) && (y < 632) );
assign R = (aW|bW)? (bW? Awins&counter[23:22]:Bwins&counter[23:22]):(white & (~black|(ball&mod1)|(wall&mod1)));
assign G = (aW|bW)? (bW? Awins&counter[23:22]:Bwins&counter[23:22]):(white & (~black|(ball&mod2)|(wall&mod2)));
assign B = (aW|bW)? (bW? Awins&~counter[23:22]:Bwins&~counter[23:22]):(white & (~black|(ball&mod3)|(wall&mod3)));

assign wall = topWall | downWall | leftWall | rightWall;
assign black = barA | barB | ball | wall | cLine;
assign white = vis;

assign check = kReg[1]^kReg[2]^kReg[3]^kReg[4]^kReg[5]^kReg[6]^kReg[7]^kReg[8]^kReg[9];

//assign PERIOD = 5000000;

//////////////////////////////////////////////////////////////////////////////////
// Design
//////////////////////////////////////////////////////////////////////////////////
// FSM
always@(posedge clk, posedge rst)
begin
	if(rst)  cState <= 0;
	else begin
		cState <= nState;
		nState <= PSCLK;
	end
end
//x
always@(posedge clk, posedge rst)
begin
    if(rst) x <= 0;
    else begin
        x <= (x < 1039)? x+1 : 0;
    end
end
// y
always@(posedge clk, posedge rst)
begin
    if(rst) y <= 0;
    else begin
        y <= (y == 665)? 0 : (x == 1039) ? y+1 : y;
    end
end
// isStop
always@(posedge clk, posedge rst)
begin
    if(rst) isStop <= 0;
    else begin
        if(sp) isStop <= ~isStop;
        else isStop <= isStop;
    end
end
// counter
always@(posedge clk, posedge rst)
begin
    if(rst) counter <= 0;
    else begin
        if(isStop) counter <= counter;
        else if(counter == PERIOD) counter <= 0;
        else counter <= counter + 1;
    end
end

/*
// ppp
always@(posedge clk, posedge rst)
begin
	if(rst) ppp <= 500000;
	else if(counter == 10) ppp <= ppp - 1;
	else ppp <= ppp;
end
*/
// PERIOD
always@(posedge clk, posedge rst)
begin
    if(rst) PERIOD <= 5000000;
    else begin
        if(counter == 5) PERIOD <= (PERIOD > 2000000)? PERIOD-20 : PERIOD;
        else PERIOD <= PERIOD;
    end
end

// timer
always@(posedge clk, posedge rst)
begin
    if(rst) timer <= 0;
    else begin
        if(timer) timer <= 0;
        else if(counter == PERIOD) timer <= 1;
        else timer <= timer;
    end
end
/*
// time2
always@(posedge clk, posedge rst)
begin
    if(rst) time2 <= 0;
    else begin
        if(time2==16) time2 <= 0;
        else if(timer) time2 <= time2+1;
        else time2 <= time2;
    end
end
*/
// kCounter
always@(posedge clk, posedge rst)
begin
	if(rst) kCounter <= 0;
	else begin
		if({cState,nState} == 2'b10) begin
			if(kCounter == 10) kCounter <= 0;
			else kCounter <= kCounter + 1;
		end else kCounter <= kCounter;
	end
end
// kReg
always@(posedge clk, posedge rst)
begin
	if(rst) kReg <= 0;
	else begin
		case({cState,nState})
			2'b10: kReg <= {PSDATA, kReg[21:1]};
			default: kReg <= kReg;
		endcase
	end
end
// kData
always@(posedge clk, posedge rst)
begin
	if(rst) kData <= 0;
	else begin
		if(kCounter == 4'd0 && check == 1'b1) begin
			if(kReg[11:1] == 11'hXX) kData <= 8'd0;
			else kData <= kReg[19:12];
		end
		else kData <= kData;
	end
end
// keyboard
always@(posedge clk, posedge rst)
begin
	if(rst) sig_f0<=0;
	else begin
		if(kData==8'hf0)sig_f0<=1;
		else if(sig_f0) begin
			case(kData)
				8'h75: up <= 1; // up
				8'h72: down <= 1; // down
                8'h6B: left <= 1; // left
                8'h74: right <= 1; // right
                8'h1d: w <= 1; // w
                8'h1b: s <= 1; // s
                8'h1c: a <= 1; // a
                8'h23: d <= 1; // d
                8'h29: sp <= 1; // space
			endcase
			sig_f0<=0;
			end
		else begin 
			sig_f0<=0;
			up<=0;
			down<=0;
            right<=0;
            left<=0;
            w<=0;
            s<=0;
            a<=0;
            d<=0;
            sp<=0;
		end
	end
end
/*
// bStepX
always@(posedge clk, posedge rst)
begin
    if(rst) bStepX <= StepXinit;
    else begin
        if(time2==16) bStepX <= (bStepX+1 < MaxSpeedX)? bStepX+1:bStepX;
        else bStepX <= bStepX;
    end
end
// bStepY
always@(posedge clk, posedge rst)
begin
    if(rst) bStepY <= StepYinit;
    else begin
        if(time2==16) bStepY <= (bStepY+1 < MaxSpeedY)? bStepY+1:bStepY;
        else bStepY <= bStepY;
    end
end
*/
// cLine
always@(posedge clk, posedge rst)
begin
    if(rst) cLine <= 0;
    else begin
        if(y > topY && y < downY && x < centerX+1 && x > centerX-1) cLine <= 1;
        else cLine <= 0;
    end
end
// topWall
always@(posedge clk, posedge rst)
begin
	if(rst) topWall <= 0;
	else begin
		if(y > topY && y < topY+wallW && x > leftX && x < rightX) topWall <= 1;
		else topWall <= 0;
	end
end
// downWall
always@(posedge clk, posedge rst)
begin
	if(rst) downWall <= 0;
	else begin
		if(y > downY-wallW && y < downY && x > leftX && x < rightX) downWall <= 1;
		else downWall <= 0;
	end
end
// leftWall
always@(posedge clk, posedge rst)
begin
	if(rst) leftWall <= 0;
	else begin
		if((y > downY-hp || y < topY+hp) && (x > leftX && x < leftX+wallW)) leftWall <= 1;
		else leftWall <= 0;
	end
end
// rightWall
always@(posedge clk, posedge rst)
begin
	if(rst) rightWall <= 0;
	else begin
		if((y > downY-hp || y < topY+hp) && (x > rightX-wallW && x < rightX)) rightWall <= 1;
		else rightWall <= 0;
	end
end

// mod1,mod2,mod3
always@(posedge clk, posedge rst)
begin
	if(rst) begin mod1 <= 1; mod2 <= 0; mod3 <= 0; end
	else begin
		if(pCenterX > rightX-radius || pCenterX < leftX+wallW+radius ||
           (pCenterY < barAy+barL+10 && pCenterY > barAy-10 && pCenterX < barAx+wallW+radius) ||
           (pCenterY < barBy+barL+10 && pCenterY > barBy-10 && pCenterX > barBx-radius) ||
		   (pCenterY < topY+wallW+radius || pCenterY > downY-wallW-radius) ) begin
			if(mod1) begin mod1 <= 0; mod2 <= 1; mod3 <=0; end
			else if(mod2) begin mod1 <= 0; mod2 <= 0; mod3 <= 1; end
			else begin mod1 <= 1; mod2 <= 0; mod3 <= 0; end
		end else begin mod1 <= mod1; mod2 <= mod2; mod3 <= mod3; end
	end
end
// ball
always@(posedge clk, posedge rst)
begin
    if(rst) ball <= 0;
    else begin
        if((x-bCenterX)*(x-bCenterX) + (y-bCenterY)*(y-bCenterY) <= radius*radius) ball <= 1;
        else ball <= 0;
    end
end
// bXd
always@(posedge clk, posedge rst)
begin
    if(rst) bXd <= 0;
    else begin
        if((pCenterY < topY+hp && pCenterY > topY && pCenterX > rightX-wallW-radius) ||
		   (pCenterY < topY+hp && pCenterY > topY && pCenterX < leftX+wallW+radius) ||
		   (pCenterY > downY-hp && pCenterY < downY && pCenterX > rightX-wallW-radius) ||
		   (pCenterY > downY-hp && pCenterY < downY && pCenterX < leftX+wallW+radius) ||
           (pCenterY < barAy+barL+10 && pCenterY > barAy-10 && pCenterX < barAx+wallW+radius) ||
           (pCenterY < barBy+barL+10 && pCenterY > barBy-10 && pCenterX > barBx-radius)) bXd <= ~bXd;
        else bXd <= bXd;
    end
end
// bYd
always@(posedge clk, posedge rst)
begin
    if(rst) bYd <= 0;
    else begin
        if(pCenterY < topY+wallW+radius || pCenterY > downY-wallW-radius)  bYd <= ~bYd;
        else bYd <= bYd;
    end
end
// bCenterX
always@(posedge clk, posedge rst)
begin
    if(rst) bCenterX <= bInitX;
    else begin
        if(timer)
            if(bXd) bCenterX <= bCenterX + bStepX;
            else bCenterX <= bCenterX - bStepX;
        else bCenterX <= bCenterX;
    end
end
// bCenterY
always@(posedge clk, posedge rst)
begin
    if(rst) bCenterY <= bInitY;
    else begin
        if(timer)
            if(bYd) bCenterY <= bCenterY + bStepY;
            else bCenterY <= bCenterY - bStepY;
        else bCenterY <= bCenterY;
    end
end
// pCenterX
assign pCenterX=(bXd)?(bCenterX + bStepX):(bCenterX - bStepX);
// pCenterY
assign pCenterY=(bYd)?(bCenterY + bStepY):(bCenterY - bStepY);
// barA
always@(posedge clk, posedge rst)
begin
    if(rst) barA <= 0;
    else begin
        if((x < barAx+barW && x > barAx) && (y < barAy+barL && y > barAy)) barA <= 1;
        else barA <= 0;
    end
end
// barB
always@(posedge clk, posedge rst)
begin
    if(rst) barB <= 0;
    else begin
        if((x < barBx+barW && x > barBx) && (y < barBy+barL && y > barBy)) barB <= 1;
        else barB <= 0;
    end
end

// barAx
always@(posedge clk, posedge rst)
begin
    if(rst) barAx <= initAX;
    else begin
        if(isStop) barAx <= barAx;
        else if(a) barAx <= (barAx-uStepX >= leftAX)? barAx-uStepX : barAx;
        else if(d) barAx <= (barAx+wallW+uStepX <= centerX)? barAx+uStepX : barAx;
        else barAx <= barAx;
    end
end
// barAy
always@(posedge clk, posedge rst)
begin
    if(rst) barAy <= initY;
    else begin
        if(isStop) barAy <= barAy;
        else if(w) barAy <= (barAy-uStepY > topY)? barAy-uStepY : barAy;
        else if(s) barAy <= (barAy+barL+uStepY < downY)? barAy+uStepY : barAy;
        else barAy <= barAy;
    end
end
// barBx
always@(posedge clk, posedge rst)
begin
    if(rst) barBx <= initBX;
    else begin
        if(isStop) barBx <= barBx;
        else if(left) barBx <= (barBx-uStepX >= centerX)? barBx-uStepX : barBx;
        else if(right) barBx <= (barBx+uStepX <= rightBX)? barBx+uStepX : barBx;
        else barBx <= barBx;
    end
end
// barBy
always@(posedge clk, posedge rst)
begin
    if(rst) barBy <= initY;
    else begin
        if(isStop) barBy <= barBy;
        else if(up) barBy <= (barBy-uStepY > topY)? barBy-uStepY : barBy;
        else if(down) barBy <= (barBy+barL+uStepY < downY)? barBy+uStepY : barBy;
        else barBy <= barBy;
    end
end
// barL
always@(posedge clk, posedge rst)
begin
    if(rst) barL <= 120;
    else begin
        if((pCenterY < barAy+barL+10 && pCenterY > barAy-10 && pCenterX < barAx+wallW+radius) ||
           (pCenterY < barBy+barL+10 && pCenterY > barBy-10 && pCenterX > barBx-radius)) barL <= (barL > 40)? barL-5:barL;
        else barL <= barL;
    end
end

// over
always@(posedge clk, posedge rst)
begin
    if(rst) begin aW <= 0; bW <= 0; end
    else begin
		if(aW == 0 && bW == 0) begin
			if(bCenterX < leftX+wallW+radius) aW <= 1;
			else if(bCenterX > rightX-radius) bW <= 1;
			else begin aW <= aW; bW <= bW; end
		end else begin aW <= aW; bW <= bW; end
    end
end

// Awins
always@(posedge clk, posedge rst)
begin
    if(rst) Awins <= 0;
    else begin
        case(y-poY)
			0: Awins <= A0[400+poX-x];
			1: Awins <= A1[400+poX-x];
			2: Awins <= A2[400+poX-x];
			3: Awins <= A3[400+poX-x];
			4: Awins <= A4[400+poX-x];
			5: Awins <= A5[400+poX-x];
			6: Awins <= A6[400+poX-x];
			7: Awins <= A7[400+poX-x];
			8: Awins <= A8[400+poX-x];
			9: Awins <= A9[400+poX-x];
			10: Awins <= A10[400+poX-x];
			11: Awins <= A11[400+poX-x];
			12: Awins <= A12[400+poX-x];
			13: Awins <= A13[400+poX-x];
			14: Awins <= A14[400+poX-x];
			15: Awins <= A15[400+poX-x];
			16: Awins <= A16[400+poX-x];
			17: Awins <= A17[400+poX-x];
			18: Awins <= A18[400+poX-x];
			19: Awins <= A19[400+poX-x];
			20: Awins <= A20[400+poX-x];
			21: Awins <= A21[400+poX-x];
			22: Awins <= A22[400+poX-x];
			23: Awins <= A23[400+poX-x];
			24: Awins <= A24[400+poX-x];
			25: Awins <= A25[400+poX-x];
			26: Awins <= A26[400+poX-x];
			27: Awins <= A27[400+poX-x];
			28: Awins <= A28[400+poX-x];
			29: Awins <= A29[400+poX-x];
			30: Awins <= A30[400+poX-x];
			31: Awins <= A31[400+poX-x];
			32: Awins <= A32[400+poX-x];
			33: Awins <= A33[400+poX-x];
			34: Awins <= A34[400+poX-x];
			35: Awins <= A35[400+poX-x];
			36: Awins <= A36[400+poX-x];
			37: Awins <= A37[400+poX-x];
			38: Awins <= A38[400+poX-x];
			39: Awins <= A39[400+poX-x];
			40: Awins <= A40[400+poX-x];
			41: Awins <= A41[400+poX-x];
			42: Awins <= A42[400+poX-x];
			43: Awins <= A43[400+poX-x];
			44: Awins <= A44[400+poX-x];
			45: Awins <= A45[400+poX-x];
			46: Awins <= A46[400+poX-x];
			47: Awins <= A47[400+poX-x];
			48: Awins <= A48[400+poX-x];
			49: Awins <= A49[400+poX-x];
			50: Awins <= A50[400+poX-x];
			51: Awins <= A51[400+poX-x];
			52: Awins <= A52[400+poX-x];
			53: Awins <= A53[400+poX-x];
			54: Awins <= A54[400+poX-x];
			55: Awins <= A55[400+poX-x];
			56: Awins <= A56[400+poX-x];
			57: Awins <= A57[400+poX-x];
			58: Awins <= A58[400+poX-x];
			59: Awins <= A59[400+poX-x];
			60: Awins <= A60[400+poX-x];
			61: Awins <= A61[400+poX-x];
			62: Awins <= A62[400+poX-x];
			63: Awins <= A63[400+poX-x];
			64: Awins <= A64[400+poX-x];
			65: Awins <= A65[400+poX-x];
			66: Awins <= A66[400+poX-x];
			67: Awins <= A67[400+poX-x];
            default: Awins <= 0;
        endcase
    end
end
// Bwins
always@(posedge clk, posedge rst)
begin
    if(rst) Bwins <= 0;
    else begin
        case(y-poY)
			0: Bwins <= B0[400+poX-x];
			1: Bwins <= B1[400+poX-x];
			2: Bwins <= B2[400+poX-x];
			3: Bwins <= B3[400+poX-x];
			4: Bwins <= B4[400+poX-x];
			5: Bwins <= B5[400+poX-x];
			6: Bwins <= B6[400+poX-x];
			7: Bwins <= B7[400+poX-x];
			8: Bwins <= B8[400+poX-x];
			9: Bwins <= B9[400+poX-x];
			10: Bwins <= B10[400+poX-x];
			11: Bwins <= B11[400+poX-x];
			12: Bwins <= B12[400+poX-x];
			13: Bwins <= B13[400+poX-x];
			14: Bwins <= B14[400+poX-x];
			15: Bwins <= B15[400+poX-x];
			16: Bwins <= B16[400+poX-x];
			17: Bwins <= B17[400+poX-x];
			18: Bwins <= B18[400+poX-x];
			19: Bwins <= B19[400+poX-x];
			20: Bwins <= B20[400+poX-x];
			21: Bwins <= B21[400+poX-x];
			22: Bwins <= B22[400+poX-x];
			23: Bwins <= B23[400+poX-x];
			24: Bwins <= B24[400+poX-x];
			25: Bwins <= B25[400+poX-x];
			26: Bwins <= B26[400+poX-x];
			27: Bwins <= B27[400+poX-x];
			28: Bwins <= B28[400+poX-x];
			29: Bwins <= B29[400+poX-x];
			30: Bwins <= B30[400+poX-x];
			31: Bwins <= B31[400+poX-x];
			32: Bwins <= B32[400+poX-x];
			33: Bwins <= B33[400+poX-x];
			34: Bwins <= B34[400+poX-x];
			35: Bwins <= B35[400+poX-x];
			36: Bwins <= B36[400+poX-x];
			37: Bwins <= B37[400+poX-x];
			38: Bwins <= B38[400+poX-x];
			39: Bwins <= B39[400+poX-x];
			40: Bwins <= B40[400+poX-x];
			41: Bwins <= B41[400+poX-x];
			42: Bwins <= B42[400+poX-x];
			43: Bwins <= B43[400+poX-x];
			44: Bwins <= B44[400+poX-x];
			45: Bwins <= B45[400+poX-x];
			46: Bwins <= B46[400+poX-x];
			47: Bwins <= B47[400+poX-x];
			48: Bwins <= B48[400+poX-x];
			49: Bwins <= B49[400+poX-x];
			50: Bwins <= B50[400+poX-x];
			51: Bwins <= B51[400+poX-x];
			52: Bwins <= B52[400+poX-x];
			53: Bwins <= B53[400+poX-x];
			54: Bwins <= B54[400+poX-x];
			55: Bwins <= B55[400+poX-x];
			56: Bwins <= B56[400+poX-x];
			57: Bwins <= B57[400+poX-x];
			58: Bwins <= B58[400+poX-x];
			59: Bwins <= B59[400+poX-x];
			60: Bwins <= B60[400+poX-x];
			61: Bwins <= B61[400+poX-x];
			62: Bwins <= B62[400+poX-x];
			63: Bwins <= B63[400+poX-x];
			64: Bwins <= B64[400+poX-x];
            default: Bwins <= 0;
        endcase
    end
end

assign A0 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign A1 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign A2 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign A3 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign A4 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign A5 = 400'b0000000000001111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000001111111111111111111100000001111111111111111111100000001111111111111111111111111111100000000000000000000000000000000001111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111100000000000000000;
assign A6 = 400'b0000000000001111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000001111111111111111111100000001111111111111111111100000001111111111111111111111111111100000000000000000000000000000000001111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111100000000000000000;
assign A7 = 400'b0000000110001111111111111111111111111111111111111111111111100000000000110000000110000000110000000110000000110001111111111111111111100000000000110000000110000000110000000110001111111111111111111100000001111111111111111111100000001111111111111111111111111111100000000000111000000111000000111001111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111100000000000000000;
assign A8 = 400'b0000011111111111111111111111111111111111111111111111111111100000000011111110011111110011111110011111110011111111111111111111111111100000000011111110011111110011111110011111111111111111111111111100000001111111111111111111100000001111111111111111111111111111100000000011111110011111110011111111111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111100000000000000000;
assign A9 = 400'b0000001111001111111111111111111111111111111111111111111111111111100001111000001111000001111000001111000001111001111111111111111111111111100001111100001111100001111100001111101111111111111111111111111101111111111111111111111111101111111111111111111111111111111111100001111100001111100001111101111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111100000000000;
assign A10 = 400'b0000001101101111111111111111111111111111111111111111111111111111100001101100001101100001101100001101100001101101111111111111111111111111100001101100001101100001101100001101101111111111111111111111111101111111111111111111111111101111111111111111111111111111111111100001101100001101100001101101111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111110000000000;
assign A11 = 400'b0000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000001111111111111111111111111101111111111111111111111111101111111111111111111111111111111111100000000000000000000000000001111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111110000000000;
assign A12 = 400'b0000000000001111111111111111111111111111111111111111111111101111100000000000000000000000000000000000000000000001111111111111111111101111100000000000000000000000000000000000001111111111111111111101111101111111111111111111101111101111111111111111111111111111101111100000000000000000000000000001111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A13 = 400'b0000011111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000001111111111111111111101111100000000000000000000000000000000000001111111111111111111101111101111111111111111111101111101111111111111111111111111111111111110000000000000000000000000001111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A14 = 400'b0001111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000001111111111111111111101111100000000000000000000000000000000000001111111111111111111101111101111111111111111111101111101111111111111111111111111111111111111100000000000000000000000001111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A15 = 400'b0001111111111111111111100000000000000000000000001111111111111111111100000000000110000000110000000110000000110001111111111111111111101111100000110000000110000000110000000110001111111111111111111101111101111111111111111111101111101111111111111111111111111111111111111100000000000010000000010001111111111111111111101111101111111111111111111100000000000000000000000000000000000000000000001111110000000000;
assign A16 = 400'b0001111111111111111111100000000000000000000000001111111111111111111100000000011111100011111100011111100011111111111111111111111111101111100011111100011111100011111100011111111111111111111111111101111101111111111111111111101111101111111111111111111111111111111111111100000000011111110011111111111111111111111111101111101111111111111111111100000000000000000000000000000000000000000000001111110000000000;
assign A17 = 400'b0001111111111111111111100000000000000000000000001111111111111111111100000000011111100011111100011111100011111101111111111111111111101111100011111100011111100011111100011111101111111111111111111101111101111111111111111111101111101111111111111111111111111111111111111100000000011111110011111111111111111111111111101111101111111111111111111100000000000000000000000000000000000000000000001111110000000000;
assign A18 = 400'b0001111111111111111111101111111111111111111111111111111111111111111111111100001111100001111100001111100001111101111111111111111111101111100001111100001111100001111100001111101111111111111111111101111101111111111111111111101111101111111111111111111111111111111111111111111100001111100001111101111111111111111111101111101111111111111111111101111111111111111111111111111111111111111111111111110000000000;
assign A19 = 400'b0001111111111111111111101111111111111111111111111111111111111111111111111100001001000001001000001001000001001001111111111111111111101111100000001000000001000000001000000001001111111111111111111101111101111111111111111111101111101111111111111111111111111111111111111111111100000001000000001001111111111111111111101111101111111111111111111101111111111111111111111111111111111111111111111111100000000000;
assign A20 = 400'b0001111111111111111111101111100000000000000000001111111111111111111101111100000000000000000000000000000000000001111111111111111111101111100000000000000000000000000000000000001111111111111111111101111101111111111111111111101111101111111111111111111111111111111111111101111100000000000000000001111111111111111111101111101111111111111111111101111110000000000000000000000000000000000000000000000000000000;
assign A21 = 400'b0001111111111111111111101111100000000000000000001111111111111111111101111100000000000000000000000000000000000001111111111111111111101111100000000000000000000000000000000000001111111111111111111101111101111111111111111111101111101111111111111111111111111111111111111101111100000000000000000001111111111111111111101111101111111111111111111101111110000000000000000000000000000000000000000000000000000000;
assign A22 = 400'b0001111111111111111111111111111111111111111111111111111111111111111101111100000000000000000000000000000000000001111111111111111111101111100000000001111111111100000000000000001111111111111111111101111101111111111111111111101111101111111111111111111111111111111111111111111111100000000000000001111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111100000000000000000;
assign A23 = 400'b0001111111111111111111111111111111111111111111111111111111111111111101111100000000000000000000000000000000000001111111111111111111101111100000000001111111111100000000000000001111111111111111111101111101111111111111111111101111101111111111111111111111111111111111111111111111100000000000000001111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111100000000000000000;
assign A24 = 400'b0001111111111111111111111111111111111111111111111111111111111111111101111100000110000000110000000110000000110001111111111111111111101111100000110001111111111100000000000110001111111111111111111101111101111111111111111111101111101111111111111111111100000001111111111111111111100000000000111001111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111100000000000000000;
assign A25 = 400'b0001111111111111111111111111111111111111111111111111111111111111111101111100011111110011111110011111110011111111111111111111111111101111100011111111111111111100000000011111111111111111111111111101111101111111111111111111101111101111111111111111111100000001111111111111111111100000000011111111111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111100000000000000000;
assign A26 = 400'b0001111111111111111111111111111111111111111111111111111111111111111101111100001111100001111100001111100001111101111111111111111111101111100001111101111111111111111100001111101111111111111111111101111101111111111111111111101111101111111111111111111101111111111111111111111111111111100001111101111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111111111100000000000;
assign A27 = 400'b0001111111111111111111111111111111111111111111111111111111111111111101111100001111100001111100001111100001111101111111111111111111101111100001111101111111111111111100001111101111111111111111111101111101111111111111111111101111101111111111111111111101111111111111111111111111111111100001111101111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111111111110000000000;
assign A28 = 400'b0001111111111111111111111111111111111111111111111111111111111111111101111100000000000000000000000000000000000001111111111111111111101111100000000001111111111111111100000000001111111111111111111101111101111111111111111111101111101111111111111111111101111111111111111111111111111111100000000001111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111111111110000000000;
assign A29 = 400'b0001111111111111111111111111111111111111111111111111111111111111111101111100000000000000000000000000000000000001111111111111111111101111100000000001111111111101111100000000001111111111111111111101111101111111111111111111101111101111111111111111111101111101111111111111111111101111100000000001111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A30 = 400'b0001111111111111111111111111111111111111111111111111111111111111111101111100000000000000000000000000000000000001111111111111111111101111100000000001111111111101111100000000001111111111111111111101111101111111111111111111101111101111111111111111111101111101111111111111111111101111100000000001111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A31 = 400'b0001111111111111111111111111111111111111111111111111111111111111111101111100000000000000000000000000000000000001111111111111111111101111101111111111111111111111111111100000001111111111111111111101111101111111111111111111101111101111111111111111111101111101111111111111111111111111111100000001111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A32 = 400'b0001111111111111111111100000000000000000000000001111111111111111111101111100000000000000000000000000000000000001111111111111111111101111101111111111111111111111111111100000001111111111111111111101111101111111111111111111101111101111111111111111111101111100001111101111111111111111111100000001111111111111111111101111100001111100000000000000000000000000000000000001111111111111111111101111110000000000;
assign A33 = 400'b0001111111111111111111100000000000000000000000001111111111111111111101111100011111100011111100011111100011111101111111111111111111101111101111111111111111111111111111100000001111111111111111111101111101111111111111111111101111101111111111111111111101111100001111101111111111111111111100000001111111111111111111101111100001111100000000000000000000000000000000000001111111111111111111101111110000000000;
assign A34 = 400'b0001111111111111111111100000000000000000000000001111111111111111111101111100011111110011111110011111110011111111111111111111111111101111101111111111111111111111111111100000001111111111111111111101111101111111111111111111101111101111111111111111111101111100001111101111111111111111111100000001111111111111111111101111100001111100000000000000000000000000000000000001111111111111111111101111110000000000;
assign A35 = 400'b0001111111111111111111101111111111111111111111111111111111111111111101111100001111000001111000001111000001111101111111111111111111101111101111111111111111111111111111111111101111111111111111111101111101111111111111111111101111101111111111111111111101111100001111111111111111111111111111111101111111111111111111101111100001111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A36 = 400'b0001111111111111111111101111111111111111111111111111111111111111111101111100001101000001101000001101000001101001111111111111111111101111101111111111111111111111111111111111101111111111111111111101111101111111111111111111101111101111111111111111111101111100001111111111111111111111111111111101111111111111111111101111100001111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A37 = 400'b0001111111111111111111101111100000000000000000001111111111111111111101111100000000000000000000000000000000000001111111111111111111101111101111111111111111111111111111101111101111111111111111111101111101111111111111111111101111101111111111111111111101111100000000001111111111111111111101111101111111111111111111101111100000000000000000000000000000000000000000000001111111111111111111101111110000000000;
assign A38 = 400'b0001111111111111111111101111100000000000000000001111111111111111111101111100000000000000000000000000000000000001111111111111111111101111101111111111111111111111111111101111101111111111111111111101111101111111111111111111101111101111111111111111111101111100000000001111111111111111111101111101111111111111111111101111100000000000000000000000000000000000000000000001111111111111111111101111110000000000;
assign A39 = 400'b0001111111111111111111101111100000000000000000001111111111111111111101111100000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101111111111111111111101111101111111111111111111101111100000000001111111111111111111111111111111111111111111111101111100111111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A40 = 400'b0001111111111111111111101111100000000000000000001111111111111111111101111100000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101111111111111111111101111101111111111111111111101111100000000001111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A41 = 400'b0001111111111111111111101111100000110000000110001111111111111111111101111100000110000000110000000110000000110000001111101111111111111111111111111111100000001111111111111111111111111111100000000001111101111111111111111111101111101111111111111111111101111100000110000001111101111111111111111111111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A42 = 400'b0001111111111111111111101111100011111100011111111111111111111111111101111100011111110011111110011111110011111110001111101111111111111111111111111111100000001111111111111111111111111111100000000001111101111111111111111111101111101111111111111111111101111100011111110001111101111111111111111111111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A43 = 400'b0001111111111111111111101111100011111100011111101111111111111111111101111100011111100011111100011111100011111100001111111111111111111111111111111111101111111111111111111111111111111111101111111111111101111111111111111111101111101111111111111111111101111100011111100001111111111111111111111111111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A44 = 400'b0001111111111111111111101111100001111100001111101111111111111111111101111100001111100001111100001111100001111100001111111111111111111111111111111111101111111111111111111111111111111111101111111111111101111111111111111111101111101111111111111111111101111100001111100001111111111111111111111111111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A45 = 400'b0001111111111111111111101111100000000000000000001111111111111111111101111100000000000000000000000000000000000000001111111111111111111111111111111111101111111111111111111111111111111111101111111111111101111111111111111111101111101111111111111111111101111100000000000001111111111111111111111111111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A46 = 400'b0001111111111111111111101111100000000000000000001111111111111111111101111100000000000000000000000000000000000000000000001111111111111111111111111111101111101111111111111111111111111111101111100000000001111111111111111111101111101111111111111111111101111100000000000000000001111111111111111111111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A47 = 400'b0001111111111111111111101111100000000000000000001111111111111111111101111100000000000000000000000000000000000000000000001111111111111111111111111111101111101111111111111111111111111111101111100000000001111111111111111111101111101111111111111111111101111100000000000000000001111111111111111111111111111111111111101111101111111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A48 = 400'b0001111111111111111111101111100000000000000000001111111111111111111101111100000000000000000000000000000000000000000000001111111111111111111111111111101111101111111111111111111111111111101111100000000001111111111111111111101111101111111111111111111101111100000000000000000001111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111101111110000000000;
assign A49 = 400'b0000111111111111111111001111100000000000000000000111111111111111111001111100000000000000000000000000000000000000000000000111111111111111111111111111001111100111111111111111111111111111001111100000000000111111111111111111001111100111111111111111111001111100000000000000000000111111111111111111111111111111111111001111100111111111111111111111111111111111111111111111111111111111111111001111110000000000;
assign A50 = 400'b0000001111100000000000001111100000110000000110000001111100000000000001111100000110000000110000000110000000110000000110000001111100000000000000000000001111100001111100000000000000000000001111100000111000001111100000000000001111100001111100000000000001111100000111000000111000001111100000000000000000000000000000001111100001111100000000000000000000000000000000000000000000000000000000001111110000000000;
assign A51 = 400'b0000001111100000000000001111100011111110011111110001111100000000000001111100011111110011111110011111110011111110011111110001111100000000000000000000001111100001111100000000000000000000001111100011111110001111100000000000001111100001111100000000000001111100011111110011111110001111100000000000000000000000000000001111100001111100000000000000000000000000000000000000000000000000000000001111110000000000;
assign A52 = 400'b0000001111111111111111111111100001111000001111000001111111111111111111111100001111000001111000001111000001111000001111000001111111111111111111111111111111100001111111111111111111111111111111100001111100001111111111111111111111100001111111111111111111111100001111100001111100001111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111110000000000;
assign A53 = 400'b0000001111111111111111111111100001111100001111100001111111111111111111111100001111100001111100001111100001111100001111100001111111111111111111111111111111100001111111111111111111111111111111100001111100001111111111111111111111100001111111111111111111111100001111100001111100001111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111110000000000;
assign A54 = 400'b0000000111111111111111111111000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000011111111111111111111111111111000000011111111111111111111111111111000000000000000011111111111111111111000000011111111111111111111000000000000000000000000011111111111111111111111111111111111111000000011111111111111011111111011111111011111111011111111011111111011111000000000000;
assign A55 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign A56 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign A57 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign A58 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign A59 = 400'b0000011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111100011111110011111110011111110011111110011111110011111110011111110000000000;
assign A60 = 400'b0000011111100011111100011111100011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110011111110000000000;
assign A61 = 400'b0000001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100000000000;
assign A62 = 400'b0000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000001001000000001000000001000000001000000101000000101000000101000000101100000101100000101100000101100000000000;
assign A63 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign A64 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign A65 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign A66 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign A67 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;


assign B0 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign B1 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign B2 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign B3 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign B4 = 400'b0000000111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000011111111111111111110000000011111111111111111110000000111111111111111111111111111110000000000000000000000000000000000111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111000000000000000000;
assign B5 = 400'b0000000111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000001111111111111111111000000000000000000000000000000000000000000011111111111111111110000000011111111111111111110000000111111111111111111111111111110000000000000000000000000000000000111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111100000000000000000;
assign B6 = 400'b0000000111111111111111111111111111111111111111111111111111111100000000000110000000110000000110000001110000001110001111111111111111111000000000001100000001100000001100000001100011111111111111111110000000011111111111111111110000000111111111111111111111111111110000000000011000000011000000011000111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111100000000000000000;
assign B7 = 400'b0000000111111111111111111111111111111111111111111111111111111100000000011111100011111100011111100111111100111111111111111111111111111000000000111111100111111100111111100111111111111111111111111110000000011111111111111111110000000111111111111111111111111111110000000001111110001111110001111111111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111100000000000000000;
assign B8 = 400'b0000000111111111111111111111111111111111111111111111111111111111111100001111000001111000001111000011111000011111001111111111111111111111111000011110000011110000011110000011110011111111111111111111111111011111111111111111111111110111111111111111111111111111111111110000111100000111100000111100111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111100000000000;
assign B9 = 400'b0000000111111111111111111111111111111111111111111111111111111111111100001111000001111000011111000011111000011111001111111111111111111111111000011111000011111000011111000011110011111111111111111111111111011111111111111111111111110111111111111111111111111111111111110000111100000111100001111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000;
assign B10 = 400'b0000000111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000011111111111111111111111111011111111111111111111111110111111111111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000;
assign B11 = 400'b0000000111111111111111111111111111111111111111111111111111111101111100000000000000000000000000000000000000000000001111111111111111111011111000000000000000000000000000000000000011111111111111111110111111011111111111111111110111110111111111111111111111111111110111110000000000000000000000000000111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111101111100000000000;
assign B12 = 400'b0000000111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000001111111111111111111011111000000000000000000000000000000000000011111111111111111110111111011111111111111111110111110111111111111111111111111111111111111100000000000000000000000000111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111101111100000000000;
assign B13 = 400'b0000001111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111011111000000000000000000000000000000000000011111111111111111110111111111111111111111111110111110111111111111111111111111111111111111110000000000000000000000000111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111011111100000000000;
assign B14 = 400'b0000000111111111111111111100000000000000000000000001111111111111111111100000000000100000000100000000100000000100001111111111111111111011111000001100000001100000001100000001100011111111111111111110111111011111111111111111110111110111111111111111111111111111111111111110000000000010000000010000111111111111111111101111111111111111111111111100000000000000000000000000000000000000000000001111100000000000;
assign B15 = 400'b0000000111111111111111111100000000000000000000000001111111111111111111100000000011111100011111100011111100111111111111111111111111111011111000111111000111111000111111000111111111111111111111111110111111011111111111111111110111110111111111111111111111111111111111111110000000001111110001111111111111111111111111101111111111111111111111111100000000000000000000000000000000000000000000001111100000000000;
assign B16 = 400'b0000000111111111111111111100111111111111111111111111111111111111111111111111000011111100011111100011111100111111111111111111111111111011111000111111000111111000111111000111111111111111111111111110111111011111111111111111110111110111111111111111111111111111111111111111111100001111110001111111111111111111111111101111111111111111111111111100111111111111111111111111111111111111111111111111100000000000;
assign B17 = 400'b0000000111111111111111111101111111111111111111111111111111111111111111111111100001111000001111000011111000011111001111111111111111111011111000011111000011111000011110000011110011111111111111111110111111011111111111111111110111110111111111111111111111111111111111111111111110000111100001111100111111111111111111101111111111111111111111111101111111111111111111111111111111111111111111111111100000000000;
assign B18 = 400'b0000000111111111111111111101111111111111111111111111111111111111111111111111100001001000001001000001011000001011001111111111111111111011111000010010000010010000010010000010010011111111111111111110111111011111111111111111110111110111111111111111111111111111111111111111111110000100100000100100111111111111111111101111111111111111111111111101111111111111111111111111111111111111111111111111100000000000;
assign B19 = 400'b0000000111111111111111111101111100000000000000000001111111111111111111101111100000000000000000000000000000000000001111111111111111111011111000000000000000000000000000000000000011111111111111111110111111011111111111111111110111110111111111111111111111111111111111111110111110000000000000000000111111111111111111101111111111111111111111111101111100000000000000000000000000000000000000000000000000000000;
assign B20 = 400'b0000000111111111111111111101111100000000000000000001111111111111111111101111100000000000000000000000000000000000001111111111111111111011111000000000000000000000000000000000000011111111111111111110111111011111111111111111110111110111111111111111111111111111111111111110111110000000000000000000111111111111111111101111111111111111111111111101111100000000000000000000000000000000000000000000000000000000;
assign B21 = 400'b0000000111111111111111111111111111111111111111111111111111111111111111101111100000000000000000000000000000000000011111111111111111111011111000000000011111111111000000000000000011111111111111111110111111111111111111111111110111110111111111111111111111111111111111111111111111100000000000000000111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111000000000000000000;
assign B22 = 400'b0000000111111111111111111111111111111111111111111111111111111111111111001111100000000000000000000000000000000000011111111111111111111011111000000000011111111111000000000000000011111111111111111110111111011111111111111111110111110111111111111111111111111111111111111111111111110000000000000000111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111100000000000000000;
assign B23 = 400'b0000000111111111111111111111111111111111111111111111111111111100000000001111100000110000000110000001110000001110001111111111111111111011111000001100011111111111000000000001100011111111111111111110111111011111111111111111110111110111111111111111111110000000111111111111111111110000000000011000111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111100000000000000000;
assign B24 = 400'b0000000111111111111111111111111111111111111111111111111111111100000000001111100011111100111111100111111100111111111111111111111111111011111000111111111111111111000000000111111111111111111111111110111111011111111111111111110111110111111111111111111110000000111111111111111111110000000011111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111100000000000000000;
assign B25 = 400'b0000000111111111111111111111111111111111111111111111111111111101111111111111100001111000001111000011111000011111001111111111111111111011111000011110011111111111111111000011110011111111111111111110111111011111111111111111110111110111111111111111111110111111111111111111111111111111110000111100111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111000000000000;
assign B26 = 400'b0000000111111111111111111111111111111111111111111111111111111101111111111111100001111000011111000011111000011111001111111111111111111011111000011111011111111111111111000011111011111111111111111110111111011111111111111111110111110111111111111111111110111111111111111111111111111111110001111100111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111100000000000;
assign B27 = 400'b0000000111111111111111111111111111111111111111111111111111111101111111111111000000000000000000000000000000000000001111111111111111111011111000000000011111111111111111000000000011111111111111111110111111011111111111111111110111110111111111111111111110111111111111111111111111111111110000000000111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111100000000000;
assign B28 = 400'b0000000111111111111111111111111111111111111111111111111111111101111100000000000000000000000000000000000000000000001111111111111111111011111000000000011111111111011111000000000011111111111111111110111111011111111111111111110111110111111111111111111110111110111111111111111111110111110000000000111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111101111100000000000;
assign B29 = 400'b0000000111111111111111111111111111111111111111111111111111111101111100000000000000000000000000000000000000000000001111111111111111111011111000000000011111111111011111000000000011111111111111111110111111011111111111111111110111110111111111111111111110111110111111111111111111110111110000000000111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111101111100000000000;
assign B30 = 400'b0000001111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111011111011111111111111111111111111111000000011111111111111111110111111111111111111111111110111110111111111111111111110111110111111111111111111111111111110000000111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111100000000000;
assign B31 = 400'b0000000111111111111111111100000000000000000000000001111111111111111111100000000000000000000000000000000000000000001111111111111111111011111011111111111111111111111111111000000011111111111111111110111111011111111111111111110111110111111111111111111110111110000111110111111111111111111110000000111111111111111111101111110001111100000000000000000000000000000000000001111111111111111111101111100000000000;
assign B32 = 400'b0000000111111111111111111100000000000000000000000001111111111111111111100000000010110000011110000011110000011111001111111111111111111011111011111111111111111111111111111000000011111111111111111110111111011111111111111111110111110111111111111111111110111110000111110111111111111111111110000000111111111111111111101111110001111100000000000000000000000000000000000001111111111111111111101111100000000000;
assign B33 = 400'b0000000111111111111111111100000000000000000000000001111111111111111111100000000011111100011111100111111100111111111111111111111111111011111011111111111111111111111111111000000011111111111111111110111111011111111111111111110111110111111111111111111110111110000111110111111111111111111110000000111111111111111111101111110001111100000000000000000000000000000000000001111111111111111111101111100000000000;
assign B34 = 400'b0000000111111111111111111101111111111111111111111111111111111111111111111111100001111000001111000011111000011111001111111111111111111011111011111111111111111111111111111111111011111111111111111110111111011111111111111111110111110111111111111111111110111110000111111111111111111111111111111110111111111111111111101111110001111111111111111111111111111111111111111111111111111111111111101111100000000000;
assign B35 = 400'b0000000111111111111111111101111111111111111111111111111111111111111111111111100001011000001011000001011000011011001111111111111111111011111011111111111111111111111111111111111011111111111111111110111111011111111111111111110111110111111111111111111110111110000111111111111111111111111111111110111111111111111111101111110001111111111111111111111111111111111111111111111111111111111111101111100000000000;
assign B36 = 400'b0000000111111111111111111101111100000000000000000001111111111111111111101111100000000000000000000000000000000000001111111111111111111011111011111111111111111111111111111011111011111111111111111110111111011111111111111111110111110111111111111111111110111110000000000111111111111111111111111110111111111111111111101111110000000000000000000000000000000000000000000001111111111111111111101111100000000000;
assign B37 = 400'b0000000111111111111111111101111100000000000000000001111111111111111111101111100000000000000000000000000000000000001111111111111111111011111011111111111111111111111111111011111011111111111111111110111111011111111111111111110111110111111111111111111110111110000000000111111111111111111110111110111111111111111111101111110000000000000000000000000000000000000000000001111111111111111111101111100000000000;
assign B38 = 400'b0000000111111111111111111111111111111111111111111111111111111111111111101111100000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111110111111011111111111111111110111110111111111111111111110111110000000000111111111111111111111111111111111111111111111101111110111111111111111111111111111111111111111111111111111111111111111111111100000000000;
assign B39 = 400'b0000000111111111111111111111111111111111111111111111111111111111111111001111100000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111110111111011111111111111111110111110111111111111111111110111110000000000111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111100000000000;
assign B40 = 400'b0000000111111111111111111111111111111111111111111111111111111100000000001111100000110000000110000000110000000110000011111111111111111111111111111111111000000011111111111111111111111111111000000000111111011111111111111111110111110111111111111111111110111110000011000000111110111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111101111100000000000;
assign B41 = 400'b0000000111111111111111111111111111111111111111111111111111111100000000001111100011111100011111100011111100111111100011111111111111111111111111111111111000000011111111111111111111111111111000000000111111011111111111111111110111110111111111111111111110111110001111110000111110111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111101111100000000000;
assign B42 = 400'b0000000111111111111111111111111111111111111111111111111111111101111111111111100011111100011111100011111100011111100011111111111111111111111111111111111011111111111111111111111111111111111011111111111111011111111111111111110111110111111111111111111110111110001111110000111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111101111100000000000;
assign B43 = 400'b0000000111111111111111111111111111111111111111111111111111111101111111111111100001111000011111000011111000011111000011111111111111111111111111111111111011111111111111111111111111111111111011111111111111011111111111111111110111110111111111111111111110111110000111110000111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111101111100000000000;
assign B44 = 400'b0000000111111111111111111111111111111111111111111111111111111101111111111111100000000000000000000000000000000000000011111111111111111111111111111111111011111111111111111111111111111111111011111111111110011111111111111111110111110111111111111111111110111110000000000000111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111101111100000000000;
assign B45 = 400'b0000000111111111111111111111111111111111111111111111111111111101111100000000000000000000000000000000000000000000000000000011111111111111111111111111111011111011111111111111111111111111111011111000000000011111111111111111110111110111111111111111111110111110000000000000000000111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111101111100000000000;
assign B46 = 400'b0000000111111111111111111111111111111111111111111111111111111101111100000000000000000000000000000000000000000000000000000011111111111111111111111111111011111011111111111111111111111111111011111000000000011111111111111111110111110111111111111111111110111110000000000000000000111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111101111100000000000;
assign B47 = 400'b0000000111111111111111111111111111111111111111111111111111111101111100000000000000000000000000000000000000000000000000000011111111111111111111111111111011111011111111111111111111111111111111111000000000011111111111111111110111110111111111111111111110111110000000000000000000111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111100000000000;
assign B48 = 400'b0000000111111111111111111111111111111111111111111111111111110001111100000000000000000000000000000000000000000000000000000001111111111111111111111111110011111001111111111111111111111111100011111000000000011111111111111111100111110011111111111111111100111110000000000000000000011111111111111111111111111111111111001111110111111111111111111111111111111111111111111111111111111111111110001111100000000000;
assign B49 = 400'b0000000001111110000000000000000000000000000000000000000000000001111100010110100010110100011111100011111000011111000011111000011111000000000000000000000011111000011111000000000000000000000011111000111110000111111000000000000111110000111110000000000000111110001011010001011010000111110000000000000000000000000000001111110001111100000000000000000000000000000000000000000000000000000000001111100000000000;
assign B50 = 400'b0000000001111110000000000000000000000000000000000000000000000001111100011111100011111100011111100011111100111111100111111100011111000000000000000000000011111000011111000000000000000000000011111001111111000111111000000000000111110000111110000000000000111110001111110001111110000111110000000000000000000000000000001111110001111100000000000000000000000000000000000000000000000000000000001111100000000000;
assign B51 = 400'b0000000001111111111111111111111111111111111111111111111111111111111100001111000001111000001111000011111000011111000011111000011111111111111111111111111111111000011111111111111111111111111111111000111110000111111111111111111111110000111111111111111111111110000111100000111100000111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111100000000000;
assign B52 = 400'b0000000001111111111111111111111111111111111111111111111111111111111100001011000001011000001011000011011000011011000011011000011111111111111111111111111111111000011111111111111111111111111111111000110110000111111111111111111111110000111111111111111111111110000111100000101100000111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111100000000000;
assign B53 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign B54 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign B55 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign B56 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign B57 = 400'b0000000000010000000010000000010000000110000000110000000110000000110000000110000000110000000110000000100000000100000000100000000100000001100000001100000001100000001100000001100000001100000001100000001000000001000000001000000001000000011000000011000000011000000011000000011000000011000000011000000010000000010000000010000000010000000110000000110000000110000000110000000110000000110000000110000000000000;
assign B58 = 400'b0000000011111110011111110011111110011111110011111100011111100011111100011111100011111100011111100011111100111111100111111100111111100111111100111111000111111000111111000111111000111111000111111000111111001111111001111111001111111001111111001111110001111110001111110001111110001111110001111110001111110011111110011111110011111110011111110011111100011111100011111100011111100011111100011111100000000000;
assign B59 = 400'b0000000001111110011111110011111110011111100011111100011111100011111100011111100011111100011111100011111100011111100111111100111111100111111000111111000111111000111111000111111000111111000111111000111111000111111001111111001111111001111110001111110001111110001111110001111110001111110001111110001111110001111110011111110011111110011111100011111100011111100011111100011111100011111100011111100000000000;
assign B60 = 400'b0000000001111100001111100001111100001111100001111100001111100001111100001111100011111100011111000011111000011111000011111000011111000011111000011111000011111000011111000011111000111111000111110000111110000111110000111110000111110000111110000111110000111110000111110000111110001111110001111100001111100001111100001111100001111100001111100001111100001111100001111100001111100011111100011111000000000000;
assign B61 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign B62 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign B63 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign B64 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;


endmodule
