`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    21:11:02 01/03/2017
// Design Name:
// Module Name:    Frogger
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module Frogger(
    input rst,
    input clk,
    input PSCLK,
    input PSDATA,
	 input START,
    output red,
    output green,
    output blue,
    output hsync,
    output vsync
);

reg [20:0] x,y;


//VGA
parameter LeftX = 104,RightX =904,TopY = 24,DownY = 587;

parameter End_Lx =  124,End_Rx =  324,End_Ty = 44,End_Dy =104;
parameter FB_Lx = LeftX,FB_Rx=RightX,FB_Ty=24,FB_Dy=104;
parameter SB_Lx = LeftX ,SB_Rx=RightX,SB_Ty=105,SB_Dy=266,SB_My=186; // white line 1 pixel
parameter TB_Lx = LeftX , TB_Rx=RightX,TB_Ty=267,TB_Dy=347;
parameter B4_Lx = LeftX ,B4_Rx=RightX,B4_Ty=348,B4_Dy=428;
parameter B5_Lx = LeftX ,B5_Rx=RightX,B5_Ty=429,B5_Dy=509;
parameter B6_Lx = LeftX ,B6_Rx=RightX,B6_Ty=510,B6_Dy=590;

reg [10:0]L1_Rx,L2_Rx,L3_Rx,L4_Rx,L5_Rx,L6_Rx,L7_Rx;
parameter step_v=81,step_h=10;

reg up,down,left,right;

reg[10:0] Frog_Rx,Frog_Ty;

reg [10:0] YC1_Rx,YC2_Rx,WT_Rx,RC1_Rx,RC2_Rx;

reg r_red,r_green,r_blue;

reg End_s,FB_s;

assign vis = (x>=LeftX) && (x<=RightX) && (y>=TopY) && (y<=DownY);
reg gameover;
reg super;

reg start;

reg over,success;




assign red = vis?(over?(success?super:gameover):r_red):0;
assign green = vis?(over?(success?super:gameover):r_green):0;
assign blue = vis?(over?(success?super:gameover):r_blue):0;

assign hsync = ~( (x >= 919) && (x < 1039) );
assign vsync = ~( (y >= 659) && (y < 665) );



parameter PERIOD=50000000;

reg [30:0] count;
reg timer;
parameter poY=TopY+200;
parameter poX=LeftX+200;
//super
wire [400:0]  su0, su1, su2, su3, su4, su5, su6, su7, su8, su9, su10, su11, su12, su13, su14, su15, su16, su17, su18, su19, su20, su21, su22, su23, su24, su25, su26, su27, su28, su29, su30, su31, su32, su33, su34, su35, su36, su37, su38, su39, su40, su41, su42, su43, su44, su45, su46, su47, su48, su49, su50, su51, su52, su53, su54, su55, su56, su57, su58, su59, su60, su61, su62, su63, su64, su65, su66, su67, su68, su69, su70, su71, su72, su73, su74, su75, su76, su77, su78, su79, su80, su81, su82, su83, su84, su85, su86, su87, su88, su89, su90, su91, su92, su93, su94, su95, su96, su97, su98, su99, su100, su101, su102, su103, su104, su105, su106, su107, su108, su109, su110, su111, su112, su113, su114, su115, su116, su117, su118, su119, su120, su121, su122, su123, su124, su125, su126, su127, su128, su129, su130, su131, su132, su133, su134, su135, su136, su137, su138, su139, su140, su141, su142, su143, su144, su145, su146, su147, su148, su149, su150, su151, su152, su153, su154, su155, su156, su157, su158, su159, su160, su161, su162, su163, su164, su165, su166, su167, su168, su169, su170, su171, su172, su173, su174, su175, su176, su177, su178, su179, su180, su181, su182, su183, su184, su185, su186, su187, su188, su189, su190, su191, su192, su193, su194, su195, su196, su197, su198, su199, su200, su201, su202, su203, su204, su205, su206, su207, su208, su209, su210, su211, su212, su213, su214, su215, su216, su217, su218, su219, su220, su221, su222, su223, su224, su225, su226, su227, su228, su229, su230, su231, su232, su233, su234, su235, su236, su237, su238, su239, su240, su241, su242, su243, su244, su245, su246, su247, su248, su249, su250, su251, su252;
assign su0 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su1 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su2 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su3 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su4 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su5 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su6 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su7 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su8 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su9 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su10 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su11 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su12 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su13 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su14 = 400'b0000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000;
assign su15 = 400'b0000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000;
assign su16 = 400'b0000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000;
assign su17 = 400'b0000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000;
assign su18 = 400'b0000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000;
assign su19 = 400'b0000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000;
assign su20 = 400'b0000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000;
assign su21 = 400'b0000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000;
assign su22 = 400'b0000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000;
assign su23 = 400'b0000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000;
assign su24 = 400'b0000000000000000000000000000000000000000001110000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000011100000000000000000000000000000000000000000;
assign su25 = 400'b0000000000000000000000000000000000000000000011100000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000001000000000001111000000000000000000000000000000000000000000;
assign su26 = 400'b0000000000000000000000000000000000000000000001110000011111111111111111111111100000000000000100001111111111111111111111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111100001000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000000111100000000000000000000000000000000000000000000;
assign su27 = 400'b0000000000000000000000000000000000000000000000111100001111111111111111111111000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000001110000000000000000000000000000000000000000000000;
assign su28 = 400'b0000000000000000000000000000000000000000000000001110001111111111111111111111000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000011100000000000000000000000000000000000000000000000;
assign su29 = 400'b0000000000000000000000000000000000000000000000000011101111111111111111111111000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100001110000000000000000000000000000000000000000000000000;
assign su30 = 400'b0000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000001111111111111111111111100000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100111100000000000000000000000000000000000000000000000000;
assign su31 = 400'b0000000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000001111111111111111111111100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111101110000000000000000000000000000000000000000000000000000;
assign su32 = 400'b0000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000001111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000;
assign su33 = 400'b0000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000001111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000000;
assign su34 = 400'b0000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000001111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su35 = 400'b0000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000001111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su36 = 400'b0000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000001111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su37 = 400'b0000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000001111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su38 = 400'b0000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000001111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su39 = 400'b0000000000000000000000000000000000000000000000000000001111111111111111111111101100000000000110001111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su40 = 400'b0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su41 = 400'b0000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su42 = 400'b0000000000000000000000000000000000000000000000000000000110101111111111111111111111111111111111111111111111110110011011000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su43 = 400'b0000000000000000000000000000000000000000000000000000000000100000111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su44 = 400'b0000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111110000000000001000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su45 = 400'b0000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su46 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000100000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su47 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su48 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su49 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000001101111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su50 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000000111001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su51 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000011110001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su52 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000000111000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su53 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000011110000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su54 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000000000111000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su55 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111111111110000000000000000000000000000000000111111111111111111111111100000000000000001100000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su56 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000001011111111111111111111111100000000000000000000000000010111111111111111111111110000000000000000000000000000000000111111111111111111111111000000000000001111000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su57 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000100000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su58 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000;
assign su59 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000;
assign su60 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000;
assign su61 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111011100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000;
assign su62 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111001111000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000;
assign su63 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000110111111111111111110000011100000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000001111111111100111111110011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000;
assign su64 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su65 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su66 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su67 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su68 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su69 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su70 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su71 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su72 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su73 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su74 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su75 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su76 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su77 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su78 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su79 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000000111100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su80 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su81 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su82 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su83 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su84 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su85 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su86 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su87 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su88 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su89 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su90 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su91 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su92 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su93 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su94 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su95 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su96 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su97 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su98 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su99 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su100 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su101 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su102 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su103 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su104 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su105 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su106 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su107 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su108 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su109 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su110 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su111 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su112 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su113 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su114 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su115 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su116 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su117 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su118 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su119 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su120 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su121 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su122 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111111000000000011111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su123 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111111000000000011111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su124 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111100000000111111110010000011111111111111111111111111111111111111111111111111111111111111111111110000001111111000000000011111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su125 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su126 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su127 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su128 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su129 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su130 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su131 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su132 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su133 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su134 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su135 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su136 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su137 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su138 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su139 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su140 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su141 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su142 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su143 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su144 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su145 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su146 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su147 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su148 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su149 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su150 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su151 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su152 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su153 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su154 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su155 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su156 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su157 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111100000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su158 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111100000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su159 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111100000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su160 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000010000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100010000000000000010000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su161 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su162 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su163 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su164 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su165 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su166 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su167 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su168 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su169 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su170 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111110000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su171 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111100000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su172 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su173 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su174 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su175 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su176 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su177 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su178 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su179 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su180 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su181 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su182 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su183 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su184 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su185 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su186 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su187 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000011001110000111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su188 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su189 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su190 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su191 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su192 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su193 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su194 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su195 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su196 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su197 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su198 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000111101111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su199 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000001110001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su200 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000111000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su201 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000001110000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su202 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000111000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su203 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000011110000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su204 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000001111111111110000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su205 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000001111111111110000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su206 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000001111111111110000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su207 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000001111111111110000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su208 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000001111111111110000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su209 = 400'b0000000000000000000000000000000000000000000111111111111111111111110010000011111111111110000000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su210 = 400'b0000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su211 = 400'b0000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su212 = 400'b0000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000011111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su213 = 400'b0000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000011111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su214 = 400'b0000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000011111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su215 = 400'b0000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000011111111111111111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su216 = 400'b0000000000000000000000000000000000000000000111111111111111111111111111111111100000000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su217 = 400'b0000000000000000000000000000000000000000000111111111111111111111111111111111101000000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su218 = 400'b0000000000000000000000000000000000000000000111111111111111111111111111111111100000000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su219 = 400'b0000000000000000000000000000000000000000000111111111111111111111111111111111110001000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su220 = 400'b0000000000000000000000000000000000000000000111111111111111111111111111111111100000000011111111111111111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000;
assign su221 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su222 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su223 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000001011111111111111111111111000000000000000000000000000000000000000000000;
assign su224 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su225 = 400'b0000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000;
assign su226 = 400'b0000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000;
assign su227 = 400'b0000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000;
assign su228 = 400'b0000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000;
assign su229 = 400'b0000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000;
assign su230 = 400'b0000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000;
assign su231 = 400'b0000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000;
assign su232 = 400'b0000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000;
assign su233 = 400'b0000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000;
assign su234 = 400'b0000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000;
assign su235 = 400'b0000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000;
assign su236 = 400'b0000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000;
assign su237 = 400'b0000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000;
assign su238 = 400'b0000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000;
assign su239 = 400'b0000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000;
assign su240 = 400'b0000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000;
assign su241 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su242 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su243 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su244 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su245 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su246 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su247 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su248 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su249 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su250 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su251 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su252 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign su253 = 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

always@(posedge clk , posedge rst)
begin
	if(rst) super<=0;
	else begin
		case(y-poY)
			0: super <= su0[400+poX-x];
1: super <= su1[400+poX-x];
2: super <= su2[400+poX-x];
3: super <= su3[400+poX-x];
4: super <= su4[400+poX-x];
5: super <= su5[400+poX-x];
6: super <= su6[400+poX-x];
7: super <= su7[400+poX-x];
8: super <= su8[400+poX-x];
9: super <= su9[400+poX-x];
10: super <= su10[400+poX-x];
11: super <= su11[400+poX-x];
12: super <= su12[400+poX-x];
13: super <= su13[400+poX-x];
14: super <= su14[400+poX-x];
15: super <= su15[400+poX-x];
16: super <= su16[400+poX-x];
17: super <= su17[400+poX-x];
18: super <= su18[400+poX-x];
19: super <= su19[400+poX-x];
20: super <= su20[400+poX-x];
21: super <= su21[400+poX-x];
22: super <= su22[400+poX-x];
23: super <= su23[400+poX-x];
24: super <= su24[400+poX-x];
25: super <= su25[400+poX-x];
26: super <= su26[400+poX-x];
27: super <= su27[400+poX-x];
28: super <= su28[400+poX-x];
29: super <= su29[400+poX-x];
30: super <= su30[400+poX-x];
31: super <= su31[400+poX-x];
32: super <= su32[400+poX-x];
33: super <= su33[400+poX-x];
34: super <= su34[400+poX-x];
35: super <= su35[400+poX-x];
36: super <= su36[400+poX-x];
37: super <= su37[400+poX-x];
38: super <= su38[400+poX-x];
39: super <= su39[400+poX-x];
40: super <= su40[400+poX-x];
41: super <= su41[400+poX-x];
42: super <= su42[400+poX-x];
43: super <= su43[400+poX-x];
44: super <= su44[400+poX-x];
45: super <= su45[400+poX-x];
46: super <= su46[400+poX-x];
47: super <= su47[400+poX-x];
48: super <= su48[400+poX-x];
49: super <= su49[400+poX-x];
50: super <= su50[400+poX-x];
51: super <= su51[400+poX-x];
52: super <= su52[400+poX-x];
53: super <= su53[400+poX-x];
54: super <= su54[400+poX-x];
55: super <= su55[400+poX-x];
56: super <= su56[400+poX-x];
57: super <= su57[400+poX-x];
58: super <= su58[400+poX-x];
59: super <= su59[400+poX-x];
60: super <= su60[400+poX-x];
61: super <= su61[400+poX-x];
62: super <= su62[400+poX-x];
63: super <= su63[400+poX-x];
64: super <= su64[400+poX-x];
65: super <= su65[400+poX-x];
66: super <= su66[400+poX-x];
67: super <= su67[400+poX-x];
68: super <= su68[400+poX-x];
69: super <= su69[400+poX-x];
70: super <= su70[400+poX-x];
71: super <= su71[400+poX-x];
72: super <= su72[400+poX-x];
73: super <= su73[400+poX-x];
74: super <= su74[400+poX-x];
75: super <= su75[400+poX-x];
76: super <= su76[400+poX-x];
77: super <= su77[400+poX-x];
78: super <= su78[400+poX-x];
79: super <= su79[400+poX-x];
80: super <= su80[400+poX-x];
81: super <= su81[400+poX-x];
82: super <= su82[400+poX-x];
83: super <= su83[400+poX-x];
84: super <= su84[400+poX-x];
85: super <= su85[400+poX-x];
86: super <= su86[400+poX-x];
87: super <= su87[400+poX-x];
88: super <= su88[400+poX-x];
89: super <= su89[400+poX-x];
90: super <= su90[400+poX-x];
91: super <= su91[400+poX-x];
92: super <= su92[400+poX-x];
93: super <= su93[400+poX-x];
94: super <= su94[400+poX-x];
95: super <= su95[400+poX-x];
96: super <= su96[400+poX-x];
97: super <= su97[400+poX-x];
98: super <= su98[400+poX-x];
99: super <= su99[400+poX-x];
100: super <= su100[400+poX-x];
101: super <= su101[400+poX-x];
102: super <= su102[400+poX-x];
103: super <= su103[400+poX-x];
104: super <= su104[400+poX-x];
105: super <= su105[400+poX-x];
106: super <= su106[400+poX-x];
107: super <= su107[400+poX-x];
108: super <= su108[400+poX-x];
109: super <= su109[400+poX-x];
110: super <= su110[400+poX-x];
111: super <= su111[400+poX-x];
112: super <= su112[400+poX-x];
113: super <= su113[400+poX-x];
114: super <= su114[400+poX-x];
115: super <= su115[400+poX-x];
116: super <= su116[400+poX-x];
117: super <= su117[400+poX-x];
118: super <= su118[400+poX-x];
119: super <= su119[400+poX-x];
120: super <= su120[400+poX-x];
121: super <= su121[400+poX-x];
122: super <= su122[400+poX-x];
123: super <= su123[400+poX-x];
124: super <= su124[400+poX-x];
125: super <= su125[400+poX-x];
126: super <= su126[400+poX-x];
127: super <= su127[400+poX-x];
128: super <= su128[400+poX-x];
129: super <= su129[400+poX-x];
130: super <= su130[400+poX-x];
131: super <= su131[400+poX-x];
132: super <= su132[400+poX-x];
133: super <= su133[400+poX-x];
134: super <= su134[400+poX-x];
135: super <= su135[400+poX-x];
136: super <= su136[400+poX-x];
137: super <= su137[400+poX-x];
138: super <= su138[400+poX-x];
139: super <= su139[400+poX-x];
140: super <= su140[400+poX-x];
141: super <= su141[400+poX-x];
142: super <= su142[400+poX-x];
143: super <= su143[400+poX-x];
144: super <= su144[400+poX-x];
145: super <= su145[400+poX-x];
146: super <= su146[400+poX-x];
147: super <= su147[400+poX-x];
148: super <= su148[400+poX-x];
149: super <= su149[400+poX-x];
150: super <= su150[400+poX-x];
151: super <= su151[400+poX-x];
152: super <= su152[400+poX-x];
153: super <= su153[400+poX-x];
154: super <= su154[400+poX-x];
155: super <= su155[400+poX-x];
156: super <= su156[400+poX-x];
157: super <= su157[400+poX-x];
158: super <= su158[400+poX-x];
159: super <= su159[400+poX-x];
160: super <= su160[400+poX-x];
161: super <= su161[400+poX-x];
162: super <= su162[400+poX-x];
163: super <= su163[400+poX-x];
164: super <= su164[400+poX-x];
165: super <= su165[400+poX-x];
166: super <= su166[400+poX-x];
167: super <= su167[400+poX-x];
168: super <= su168[400+poX-x];
169: super <= su169[400+poX-x];
170: super <= su170[400+poX-x];
171: super <= su171[400+poX-x];
172: super <= su172[400+poX-x];
173: super <= su173[400+poX-x];
174: super <= su174[400+poX-x];
175: super <= su175[400+poX-x];
176: super <= su176[400+poX-x];
177: super <= su177[400+poX-x];
178: super <= su178[400+poX-x];
179: super <= su179[400+poX-x];
180: super <= su180[400+poX-x];
181: super <= su181[400+poX-x];
182: super <= su182[400+poX-x];
183: super <= su183[400+poX-x];
184: super <= su184[400+poX-x];
185: super <= su185[400+poX-x];
186: super <= su186[400+poX-x];
187: super <= su187[400+poX-x];
188: super <= su188[400+poX-x];
189: super <= su189[400+poX-x];
190: super <= su190[400+poX-x];
191: super <= su191[400+poX-x];
192: super <= su192[400+poX-x];
193: super <= su193[400+poX-x];
194: super <= su194[400+poX-x];
195: super <= su195[400+poX-x];
196: super <= su196[400+poX-x];
197: super <= su197[400+poX-x];
198: super <= su198[400+poX-x];
199: super <= su199[400+poX-x];
200: super <= su200[400+poX-x];
201: super <= su201[400+poX-x];
202: super <= su202[400+poX-x];
203: super <= su203[400+poX-x];
204: super <= su204[400+poX-x];
205: super <= su205[400+poX-x];
206: super <= su206[400+poX-x];
207: super <= su207[400+poX-x];
208: super <= su208[400+poX-x];
209: super <= su209[400+poX-x];
210: super <= su210[400+poX-x];
211: super <= su211[400+poX-x];
212: super <= su212[400+poX-x];
213: super <= su213[400+poX-x];
214: super <= su214[400+poX-x];
215: super <= su215[400+poX-x];
216: super <= su216[400+poX-x];
217: super <= su217[400+poX-x];
218: super <= su218[400+poX-x];
219: super <= su219[400+poX-x];
220: super <= su220[400+poX-x];
221: super <= su221[400+poX-x];
222: super <= su222[400+poX-x];
223: super <= su223[400+poX-x];
224: super <= su224[400+poX-x];
225: super <= su225[400+poX-x];
226: super <= su226[400+poX-x];
227: super <= su227[400+poX-x];
228: super <= su228[400+poX-x];
229: super <= su229[400+poX-x];
230: super <= su230[400+poX-x];
231: super <= su231[400+poX-x];
232: super <= su232[400+poX-x];
233: super <= su233[400+poX-x];
234: super <= su234[400+poX-x];
235: super <= su235[400+poX-x];
236: super <= su236[400+poX-x];
237: super <= su237[400+poX-x];
238: super <= su238[400+poX-x];
239: super <= su239[400+poX-x];
240: super <= su240[400+poX-x];
241: super <= su241[400+poX-x];
242: super <= su242[400+poX-x];
243: super <= su243[400+poX-x];
244: super <= su244[400+poX-x];
245: super <= su245[400+poX-x];
246: super <= su246[400+poX-x];
247: super <= su247[400+poX-x];
248: super <= su248[400+poX-x];
249: super <= su249[400+poX-x];
250: super <= su250[400+poX-x];
251: super <= su251[400+poX-x];
252: super <= su252[400+poX-x];
default: super<=0;
		endcase
	end
end

//gameover
wire [399:0]  go0, go1, go2, go3, go4, go5, go6, go7, go8, go9, go10, go11, go12, go13, go14, go15, go16, go17, go18, go19, go20, go21, go22, go23, go24, go25, go26, go27, go28, go29, go30, go31, go32, go33, go34, go35, go36, go37, go38, go39, go40, go41, go42, go43, go44, go45, go46, go47, go48, go49, go50, go51, go52, go53, go54, go55, go56, go57, go58, go59, go60, go61, go62, go63, go64, go65, go66, go67, go68, go69, go70, go71, go72, go73, go74, go75, go76, go77, go78, go79, go80, go81, go82, go83, go84, go85, go86, go87, go88, go89, go90, go91, go92, go93, go94, go95, go96, go97, go98, go99, go100, go101, go102, go103, go104, go105, go106, go107, go108, go109, go110, go111, go112, go113, go114, go115, go116, go117, go118, go119, go120, go121, go122, go123, go124, go125, go126, go127, go128, go129, go130, go131, go132, go133, go134;
assign go0 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go1 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go2 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go3 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go4 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go5 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go6 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go7 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go8 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go9 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go10 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go11 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go12 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go13 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go14 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go15 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go16 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go17 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go18 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go19 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go20 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go21 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go22 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go23 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go24 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go25 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go26 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go27 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go28 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go29 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go30 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go31 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go32 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go33 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go34 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go35 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go36 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go37 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go38 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go39 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go40 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go41 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000001111110000011111100000000000000000000000000000000000000000000000011111100000111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go42 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000001111111100111111100000000000000000000000000000000000000000000000011111110011111111000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go43 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go44 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go45 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go46 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go47 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go48 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000001111111100111111100000000000000000000000000000000000000000000000011111110011111111000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go49 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000001111110000011111100000000000000000000000000000000000000000000000011111100000111111000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go50 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go51 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go52 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go53 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go54 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go55 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go56 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go57 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go58 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go59 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go60 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go61 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go62 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go63 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go64 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go65 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go66 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go67 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go68 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go69 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go70 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go71 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go72 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go73 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go74 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go75 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000011111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go76 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000011111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go77 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000011111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go78 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000011111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go79 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000011111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go80 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000011111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go81 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000011111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go82 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go83 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go84 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go85 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go86 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go87 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go88 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go89 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go90 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go91 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go92 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go93 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go94 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go95 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111000000000100011111111011111111111111111111111111110000000000000000000001111111111111111110000000000000111111100000011111111100000001110000000000000000000000111000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go96 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111100111111111111001111111110011111111001111111111111111111110011100000001111111111111111111111111111111100011111111000111111100000001111111100000001110000000111111111111111111000000011111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go97 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111100000011110000001111111110000001111000000111111111111100000011100000001111111111111111111111111111000000011111111100000011100000001111111100000001110000000111111111111111111000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go98 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111100000011110000001111111110000001111000000111111111111100000011100000001111111111111111111111111111000000011111111100000011100000001111111100000001110000000111111111111111111000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go99 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111100000011110000001111111110000001111000000000011111000000000011100000001111111111111111111111111111000000011111111100000011100000001111111100000001110000000111111111111111111000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go100 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111110000001111111110000001111000000000011111000000000011100000001111111111111111111111111111000000011111111100000011100000001111111100000001110000000111111111111111111000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go101 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111110000001111111110000001111000000000000000000000000011100000001111111111111111111111111111000000011111111100000011100000001111111100000001110000000111111111111111111000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go102 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111110000001111111110000001111000000111110011111100000011100000001111111111111111111111111111000000011111111100000011100000001111111100000001110000000111111111111111111000000011111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go103 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111000000000011110000001111111110000001111000000111110011111100000011100000000000000000011111111111111111000000011111111100000011100000001111111100000001110000000000000000001111111000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go104 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111100000011110000001111111110000001111000000111111111111100000011100000001111111111111111111111111111000000011111111100000011111110001111111100011111110000000111111111111111111000000011111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go105 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111100000011110000000000000000000001111000000111111111111100000011100000001111111111111111111111111111000000011111111100000011111110000000000000011111110000000111111111111111111000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go106 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111100000011110000001111111110000001111000000111111111111100000011100000001111111111111111111111111111000000011111111100000011111110000000000000011111110000000111111111111111111000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go107 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111100000011110000001111111110000001111000000111111111111100000011100000001111111111111111111111111111000000011111111100000011111110000000000000011111110000000111111111111111111000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go108 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111100000011110000001111111110000001111000000111111111111100000011100000001111111111111111111111111111000000011111111100000011111111111000000111111111110000000111111111111111111000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go109 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111100000011110000001111111110000001111000000111111111111100000011100000001111111111111111111111111111000000011111111100000011111111111000000111111111110000000111111111111111111000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go110 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111100111111110000001111111110000001111000000111111111111100000011100000001111111111111111111111111111111100011111111000111111111111111000000111111111110000000111111111111111111000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go111 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111110000001111111110000001111000000111111111111100000011100000000000000000000001111111111111111100000000000000111111111111111000000111111111110000000000000000000000111000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go112 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go113 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go114 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go115 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go116 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go117 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go118 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go119 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go120 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go121 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go122 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go123 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go124 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go125 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go126 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go127 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go128 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go129 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go130 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go131 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go132 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go133 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
assign go134 = 400'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;


always@(posedge clk or posedge rst)
begin
    if(rst) gameover<=0;
    else 
		case(y-poY)
			0: gameover <= go0[400+poX-x];
1: gameover <= go1[400+poX-x];
2: gameover <= go2[400+poX-x];
3: gameover <= go3[400+poX-x];
4: gameover <= go4[400+poX-x];
5: gameover <= go5[400+poX-x];
6: gameover <= go6[400+poX-x];
7: gameover <= go7[400+poX-x];
8: gameover <= go8[400+poX-x];
9: gameover <= go9[400+poX-x];
10: gameover <= go10[400+poX-x];
11: gameover <= go11[400+poX-x];
12: gameover <= go12[400+poX-x];
13: gameover <= go13[400+poX-x];
14: gameover <= go14[400+poX-x];
15: gameover <= go15[400+poX-x];
16: gameover <= go16[400+poX-x];
17: gameover <= go17[400+poX-x];
18: gameover <= go18[400+poX-x];
19: gameover <= go19[400+poX-x];
20: gameover <= go20[400+poX-x];
21: gameover <= go21[400+poX-x];
22: gameover <= go22[400+poX-x];
23: gameover <= go23[400+poX-x];
24: gameover <= go24[400+poX-x];
25: gameover <= go25[400+poX-x];
26: gameover <= go26[400+poX-x];
27: gameover <= go27[400+poX-x];
28: gameover <= go28[400+poX-x];
29: gameover <= go29[400+poX-x];
30: gameover <= go30[400+poX-x];
31: gameover <= go31[400+poX-x];
32: gameover <= go32[400+poX-x];
33: gameover <= go33[400+poX-x];
34: gameover <= go34[400+poX-x];
35: gameover <= go35[400+poX-x];
36: gameover <= go36[400+poX-x];
37: gameover <= go37[400+poX-x];
38: gameover <= go38[400+poX-x];
39: gameover <= go39[400+poX-x];
40: gameover <= go40[400+poX-x];
41: gameover <= go41[400+poX-x];
42: gameover <= go42[400+poX-x];
43: gameover <= go43[400+poX-x];
44: gameover <= go44[400+poX-x];
45: gameover <= go45[400+poX-x];
46: gameover <= go46[400+poX-x];
47: gameover <= go47[400+poX-x];
48: gameover <= go48[400+poX-x];
49: gameover <= go49[400+poX-x];
50: gameover <= go50[400+poX-x];
51: gameover <= go51[400+poX-x];
52: gameover <= go52[400+poX-x];
53: gameover <= go53[400+poX-x];
54: gameover <= go54[400+poX-x];
55: gameover <= go55[400+poX-x];
56: gameover <= go56[400+poX-x];
57: gameover <= go57[400+poX-x];
58: gameover <= go58[400+poX-x];
59: gameover <= go59[400+poX-x];
60: gameover <= go60[400+poX-x];
61: gameover <= go61[400+poX-x];
62: gameover <= go62[400+poX-x];
63: gameover <= go63[400+poX-x];
64: gameover <= go64[400+poX-x];
65: gameover <= go65[400+poX-x];
66: gameover <= go66[400+poX-x];
67: gameover <= go67[400+poX-x];
68: gameover <= go68[400+poX-x];
69: gameover <= go69[400+poX-x];
70: gameover <= go70[400+poX-x];
71: gameover <= go71[400+poX-x];
72: gameover <= go72[400+poX-x];
73: gameover <= go73[400+poX-x];
74: gameover <= go74[400+poX-x];
75: gameover <= go75[400+poX-x];
76: gameover <= go76[400+poX-x];
77: gameover <= go77[400+poX-x];
78: gameover <= go78[400+poX-x];
79: gameover <= go79[400+poX-x];
80: gameover <= go80[400+poX-x];
81: gameover <= go81[400+poX-x];
82: gameover <= go82[400+poX-x];
83: gameover <= go83[400+poX-x];
84: gameover <= go84[400+poX-x];
85: gameover <= go85[400+poX-x];
86: gameover <= go86[400+poX-x];
87: gameover <= go87[400+poX-x];
88: gameover <= go88[400+poX-x];
89: gameover <= go89[400+poX-x];
90: gameover <= go90[400+poX-x];
91: gameover <= go91[400+poX-x];
92: gameover <= go92[400+poX-x];
93: gameover <= go93[400+poX-x];
94: gameover <= go94[400+poX-x];
95: gameover <= go95[400+poX-x];
96: gameover <= go96[400+poX-x];
97: gameover <= go97[400+poX-x];
98: gameover <= go98[400+poX-x];
99: gameover <= go99[400+poX-x];
100: gameover <= go100[400+poX-x];
101: gameover <= go101[400+poX-x];
102: gameover <= go102[400+poX-x];
103: gameover <= go103[400+poX-x];
104: gameover <= go104[400+poX-x];
105: gameover <= go105[400+poX-x];
106: gameover <= go106[400+poX-x];
107: gameover <= go107[400+poX-x];
108: gameover <= go108[400+poX-x];
109: gameover <= go109[400+poX-x];
110: gameover <= go110[400+poX-x];
111: gameover <= go111[400+poX-x];
112: gameover <= go112[400+poX-x];
113: gameover <= go113[400+poX-x];
114: gameover <= go114[400+poX-x];
115: gameover <= go115[400+poX-x];
116: gameover <= go116[400+poX-x];
117: gameover <= go117[400+poX-x];
118: gameover <= go118[400+poX-x];
119: gameover <= go119[400+poX-x];
120: gameover <= go120[400+poX-x];
121: gameover <= go121[400+poX-x];
122: gameover <= go122[400+poX-x];
123: gameover <= go123[400+poX-x];
124: gameover <= go124[400+poX-x];
125: gameover <= go125[400+poX-x];
126: gameover <= go126[400+poX-x];
127: gameover <= go127[400+poX-x];
128: gameover <= go128[400+poX-x];
129: gameover <= go129[400+poX-x];
130: gameover <= go130[400+poX-x];
131: gameover <= go131[400+poX-x];
132: gameover <= go132[400+poX-x];
133: gameover <= go133[400+poX-x];
134: gameover <= go134[400+poX-x];
			default:gameover<=0;
		endcase
end

always@(posedge clk or posedge rst)
begin
	if(rst) start<=0;
	else if(START)start<=1;
	else start<=start;
end
//counter
always@(posedge clk or posedge rst)
begin
    if(rst) count<=0;
	 else if(!start)count<=0;
    else if(count==PERIOD) count<=0;
    else count<=count+1;
end
//timer

always@(posedge clk or posedge rst)
begin
    if(rst)timer<=0;
	 else if(!start)timer<=0;
    else if(timer) timer<=0;
    else if(count==PERIOD) timer<=1;
    else timer<=timer;
end

//gameover

always @ (posedge clk, posedge rst)
begin
    if(rst) begin
        over<=0;
		  success<=0;
    end
	 else if(!start)
	 begin
		over<=0;
		success<=0;
	 end
    else if(x>=Frog_Rx && x<=Frog_Rx+60 
				&& y>=Frog_Ty && y<=Frog_Ty+60 && !success && !over)
		begin
			
        if(x>=End_Lx && x<=End_Rx && y>=End_Ty && y<=End_Dy)
				begin 
					success<=1;
					over<=1;
				end
        else if(y<=SB_My && y>=SB_Ty)
					begin
						if(y>=(SB_My-10) || y<=(SB_Ty+10))
							;
						else if( (L1_Rx+60<=RightX && x<=L1_Rx+60 && x>=L1_Rx)||
							 (L1_Rx+60>RightX && ((x<=(L1_Rx+60-RightX+LeftX) && x>=LeftX) || (x>=L1_Rx && x<=RightX))))
							;
						else if(    (L2_Rx+60<=RightX && x<=L2_Rx+60 && x>=L2_Rx)||
							 (L2_Rx+60>RightX && ((x<=(L2_Rx+60-RightX+LeftX) && x>=LeftX) || (x>=L2_Rx && x<=RightX))))
							;
						else if(    (L3_Rx+60<=RightX && x<=L3_Rx+60 && x>=L3_Rx)||
							 (L3_Rx+60>RightX && ((x<=(L3_Rx+60-RightX+LeftX) && x>=LeftX) || (x>=L3_Rx && x<=RightX))))
							;
						else if(    (L4_Rx+60<=RightX && x<=L4_Rx+60 && x>=L4_Rx)||
							 (L4_Rx+60>RightX && ((x<=(L4_Rx+60-RightX+LeftX) && x>=LeftX) || (x>=L4_Rx && x<=RightX))))
							;
						else	over<=1; 
				  end
        else if(y<=SB_Dy && y>=SB_My) 
						begin
						if(y>=(SB_Dy-10) || y<=(SB_My+10))
							;
						else if( (L5_Rx+60<=RightX && x<=L5_Rx+60 && x>=L5_Rx)||
							 (L5_Rx+60>RightX && ((x<=(LeftX+L5_Rx+60-RightX) && x>=LeftX) || (x>=L5_Rx && x<=RightX))))
					  ;
						else if(        (L6_Rx+60<=RightX && x<=L6_Rx+60 && x>=L6_Rx)||
							 (L6_Rx+60>RightX && ((x<=(LeftX+L6_Rx+60-RightX) && x>=LeftX) || (x>=L6_Rx && x<=RightX))))
					  ;
						else if(        (L7_Rx+60<=RightX && x<=L7_Rx+60 && x>=L7_Rx)||
							 (L7_Rx+60>RightX && ((x<=(LeftX+L7_Rx+60-RightX) && x>=LeftX) || (x>=L7_Rx && x<=RightX))))
						;
						else over<=1;
				  end
			else if (y<=TB_Dy && y>=TB_Ty) 
				begin
					if(y>=(TB_Dy-10) || y<=(TB_Ty+10))
							;
					else if( (WT_Rx+120<=RightX && x<=WT_Rx+120 && x>=WT_Rx)||
						  (WT_Rx+120>RightX && ((x<=(WT_Rx+120-RightX+LeftX) && x>=LeftX) 
						  || (x>=WT_Rx && x<=RightX))))
								begin over<=1; end
				end
			else if( y<=B4_Dy && y>=B4_Ty ) 
						begin
						if(y>=(B4_Dy-10) || y<=(B4_Ty+10))
						 ;
						else if( (YC1_Rx+120<=RightX && x<=YC1_Rx+120 && x>=YC1_Rx)||
							  (YC1_Rx+120>RightX && ((x<=(LeftX+YC1_Rx+120-RightX)
							  && x>=LeftX) || (x>=YC1_Rx && x<=RightX))))
							  begin over<=1; end
						 else if((YC2_Rx+120<=RightX && x<=YC2_Rx+120 && x>=YC2_Rx)||
									(YC2_Rx+120>RightX && ((x<=(LeftX+YC2_Rx+120-RightX) && x>=LeftX) 
									|| (x>=YC2_Rx && x<=RightX))))
						 begin over<=1; end
					end
			else if( y<=B5_Dy && y>=B5_Ty ) 
					begin
						if(y>=(B5_Dy-10) || y<=(B5_Ty+10))
						;
						else if( (RC1_Rx+120<=RightX && x<=RC1_Rx+120 && x>=RC1_Rx)||
										 (RC1_Rx+120>RightX && ((x<=(RC1_Rx+120-RightX+LeftX) 
										 && x>=LeftX) || (x>=RC1_Rx && x<=RightX))))
								over<=1;
					else if( (RC2_Rx+120<=RightX && x<=RC2_Rx+120 && x>=RC2_Rx)||
										 (RC2_Rx+120>RightX && ((x<=(RC2_Rx+120-RightX+LeftX) 
										 && x>=LeftX) || (x>=RC2_Rx && x<=RightX))))
								over<=1;
					end
			end
		end


//



always @ (posedge clk, posedge rst)
begin
    if(rst) begin
        r_red<=0;
        r_green<=0;
        r_blue<=0;
    end
    else begin
		  if(over)begin
			r_red<=0;r_green<=0;r_blue<=0;
		  end
		  else if(x>=Frog_Rx && x<=Frog_Rx+60 && y>=Frog_Ty && y<=Frog_Ty+60)
		  begin
		      r_red<=1;r_green<=0;r_blue<=1;
		  end
        else if(x>=End_Lx && x<=End_Rx && y>=End_Ty && y<=End_Dy)
        begin 
				r_red<=0;  r_green<=0;  r_blue<=0;
			end
        else if(x>=FB_Lx && x<=FB_Rx && y>=FB_Ty && y<=FB_Dy)
        begin r_red<=0;  r_green<=1;  r_blue<=0;end
        else if(y<SB_My && y>=SB_Ty)begin
				if(y>=(SB_My-10) || y<=(SB_Ty+10))
					begin r_red<=0;r_green<=0; r_blue<=1;end
            else if( (L1_Rx+60<=RightX && x<=L1_Rx+60 && x>=L1_Rx)||
                (L1_Rx+60>RightX && ((x<=(L1_Rx+60-RightX+LeftX) && x>=LeftX) || (x>=L1_Rx && x<=RightX))))
            begin r_red<=0;r_green<=1;r_blue<=0; end
            else if(    (L2_Rx+60<=RightX && x<=L2_Rx+60 && x>=L2_Rx)||
                (L2_Rx+60>RightX && ((x<=(L2_Rx+60-RightX+LeftX) && x>=LeftX) || (x>=L2_Rx && x<=RightX))))
            begin r_red<=0;r_green<=1;r_blue<=0; end
            else if(    (L3_Rx+60<=RightX && x<=L3_Rx+60 && x>=L3_Rx)||
                (L3_Rx+60>RightX && ((x<=(L3_Rx+60-RightX+LeftX) && x>=LeftX) || (x>=L3_Rx && x<=RightX))))
            begin r_red<=0;r_green<=1;r_blue<=0; end
            else if(    (L4_Rx+60<=RightX && x<=L4_Rx+60 && x>=L4_Rx)||
                (L4_Rx+60>RightX && ((x<=(L4_Rx+60-RightX+LeftX) && x>=LeftX) || (x>=L4_Rx && x<=RightX))))
            begin r_red<=0;r_green<=1;r_blue<=0; end
            else begin r_red<=0;r_green<=0;r_blue<=1;end
        end
        else if(y<SB_Dy && y>=SB_My) begin
				if(y>=(SB_Dy-10) || y<=(SB_My+10))
					begin r_red<=0;r_green<=0; r_blue<=1;end
            else if( (L5_Rx+60<=RightX && x<=L5_Rx+60 && x>=L5_Rx)||
                (L5_Rx+60>RightX && ((x<=(LeftX+L5_Rx+60-RightX) && x>=LeftX) || (x>=L5_Rx && x<=RightX))))
            begin r_red<=0;r_green<=1;r_blue<=0; end
            else if(        (L6_Rx+60<=RightX && x<=L6_Rx+60 && x>=L6_Rx)||
                (L6_Rx+60>RightX && ((x<=(LeftX+L6_Rx+60-RightX) && x>=LeftX) || (x>=L6_Rx && x<=RightX))))
            begin r_red<=0;r_green<=1;r_blue<=0; end
            else if(        (L7_Rx+60<=RightX && x<=L7_Rx+60 && x>=L7_Rx)||
                (L7_Rx+60>RightX && ((x<=(LeftX+L7_Rx+60-RightX) && x>=LeftX) || (x>=L7_Rx && x<=RightX))))
            begin r_red<=0;r_green<=1;r_blue<=0; end
            else begin r_red<=0;r_green<=0;r_blue<=1;end
        end
    

else if (y<TB_Dy && y>=TB_Ty) begin
	if(y>=(TB_Dy-10) || y<=(TB_Ty+10))
			begin r_red<=0;r_green<=1;r_blue<=0; end
	else if( (WT_Rx+120<=RightX && x<=WT_Rx+120 && x>=WT_Rx)||
        (WT_Rx+120>RightX && ((x<=(WT_Rx+120-RightX+LeftX) && x>=LeftX) 
		  || (x>=WT_Rx && x<=RightX))))
            begin r_red<=1;r_green<=1;r_blue<=1; end
	else 
		begin r_red<=0;r_green<=1;r_blue<=0; end
end
else if( y<B4_Dy && y>=B4_Ty ) begin
	if(y>=(B4_Dy-10) || y<=(B4_Ty+10))
	begin r_red<=0;r_green<=0;r_blue<=0; end
	else if( (YC1_Rx+120<=RightX && x<=YC1_Rx+120 && x>=YC1_Rx)||
        (YC1_Rx+120>RightX && ((x<=(LeftX+YC1_Rx+120-RightX)
		  && x>=LeftX) || (x>=YC1_Rx && x<=RightX))))
        begin r_red<=1;r_green<=1;r_blue<=0; end
    else if((YC2_Rx+120<=RightX && x<=YC2_Rx+120 && x>=YC2_Rx)||
            (YC2_Rx+120>RightX && ((x<=(LeftX+YC2_Rx+120-RightX) && x>=LeftX) 
				|| (x>=YC2_Rx && x<=RightX))))
    begin r_red<=1;r_green<=1;r_blue<=0; end
	else begin r_red<=0;r_green<=0;r_blue<=0;end
end
else if( y<B5_Dy && y>=B5_Ty ) begin
	if(y>=(B5_Dy-10) || y<=(B5_Ty+10))
	begin r_red<=0;r_green<=0;r_blue<=0; end
	else if( (RC1_Rx+120<=RightX && x<=RC1_Rx+120 && x>=RC1_Rx)||
                (RC1_Rx+120>RightX && ((x<=(RC1_Rx+120-RightX+LeftX) 
					 && x>=LeftX) || (x>=RC1_Rx && x<=RightX))))
         begin r_red<=1;r_green<=0;r_blue<=0; end
else if( (RC2_Rx+120<=RightX && x<=RC2_Rx+120 && x>=RC2_Rx)||
                (RC2_Rx+120>RightX && ((x<=(RC2_Rx+120-RightX+LeftX) 
					 && x>=LeftX) || (x>=RC2_Rx && x<=RightX))))
         begin r_red<=1;r_green<=0;r_blue<=0; end
	else 
		begin r_red<=0;r_green<=0;r_blue<=0; end
end
else if( y<B6_Dy && y>=B6_Ty ) begin
	r_red<=0;r_green<=0;r_blue<=0;
end

else if(vis) begin
    r_red<=1;r_green<=1;r_blue<=1;
end
else begin
    r_red<=0;r_green<=0;r_blue<=0;
end
end
end


    //x
always @ (posedge clk, posedge rst)
begin
    if(rst) x <= 0;
    else begin
        x <= (x < 1039)? x+1 : 0;
    end
end

// y
always @ (posedge clk, posedge rst)
begin
    if(rst) y <= 0;
    else begin
        y <= (y == 665)? 0 : (x == 1039) ? y+1 : y;
    end
end

//Frog_x
always@(posedge clk , posedge rst)
begin
	if(rst) Frog_Rx<=824;
	  else if(!start)
	 begin
			Frog_Rx<=824;	 
	end
	else begin
		if(left) Frog_Rx<=(Frog_Rx-step_h>=LeftX)?Frog_Rx-step_h:Frog_Rx;
		else if(right) Frog_Rx<=(Frog_Rx+step_h<=RightX)?Frog_Rx+step_h:Frog_Rx;
		 else if(Frog_Ty==(SB_My+10) && timer) Frog_Rx<=Frog_Rx-8;
		 else if(Frog_Ty==(SB_Ty+10) && timer) Frog_Rx<=Frog_Rx+8;
		else Frog_Rx<=Frog_Rx;
	end
end

//Frog_y

always@(posedge clk , posedge rst)
begin
	if(rst) Frog_Ty<=520;
	  else if(!start)
	 begin
			Frog_Ty<=520;	 
	end
	else begin
		if(up) Frog_Ty<=(Frog_Ty-step_v>=TopY)?Frog_Ty-step_v:Frog_Ty;
		else if(down) Frog_Ty<=(Frog_Ty+step_v<=DownY)?Frog_Ty+step_v:Frog_Ty;
		else Frog_Ty<=Frog_Ty;
	end
end



//L1_Rx
always@(posedge clk ,posedge rst)
begin
        if(rst) L1_Rx<=220;
        else begin
            if(timer) begin
                if(L1_Rx<=RightX-8)
                    L1_Rx<=L1_Rx+8;
                else
                    L1_Rx<=L1_Rx+8-RightX+LeftX;
            end
            else L1_Rx<=L1_Rx;
        end
end

//L2_Rx
always@(posedge clk ,posedge rst)
begin
    if(rst) L2_Rx<=280;
    else begin
        if(timer) begin
            if(L2_Rx<=RightX-8)
                L2_Rx<=L2_Rx+8;
            else
                L2_Rx<=L2_Rx+8-RightX+LeftX;
        end
        else L2_Rx<=L2_Rx;
    end
end

        //L3_Rx
        always@(posedge clk ,posedge rst)
        begin
            if(rst) L3_Rx<=660;
            else begin
                if(timer) begin
                    if(L3_Rx<=RightX-8)
                        L3_Rx<=L3_Rx+8;
                    else
                        L3_Rx<=L3_Rx+8-RightX+LeftX;
                end
                else L3_Rx<=L3_Rx;
            end
    end

    //L4_Rx
always@(posedge clk ,posedge rst)
    begin
        if(rst) L4_Rx<=720;
        else begin
            if(timer) begin
                if(L4_Rx<=RightX-8)
                    L4_Rx<=L4_Rx+8;
                else
                    L4_Rx<=L4_Rx+8-RightX+LeftX;
            end
            else L4_Rx<=L4_Rx;
        end
end




//L5_Rx
always@(posedge clk ,posedge rst)
begin
    if(rst) L5_Rx<=510;
    else begin
        if(timer) begin
            if(L5_Rx>=LeftX+8)
                L5_Rx<=L5_Rx-8;
            else
                L5_Rx<=RightX+(L5_Rx-LeftX-8);
        end
        else L5_Rx<=L5_Rx;
    end
end

        //L6_Rx
always@(posedge clk ,posedge rst)
 begin
            if(rst) L6_Rx<=570;
            else begin
                if(timer) begin
                    if(L6_Rx>=LeftX+8)
                        L6_Rx<=L6_Rx-8;
                    else
                        L6_Rx<=RightX+(L6_Rx-LeftX-8);
                end
                else L6_Rx<=L6_Rx;
            end
 end

    //L7_Rx
always@(posedge clk ,posedge rst)
begin
        if(rst) L7_Rx<=630;
        else begin
            if(timer) begin
                if(L7_Rx>=LeftX+8)
                    L7_Rx<=L7_Rx-8;
                else
                    L7_Rx<=RightX+(L7_Rx-LeftX-8);
            end
            else L7_Rx<=L7_Rx;
        end
end
//WT_Rx
always@(posedge clk ,posedge rst)
    begin
        if(rst) WT_Rx<=LeftX;
        else begin
            if(timer) begin
                if(WT_Rx<=RightX-6)
                    WT_Rx<=WT_Rx+6;
                else
                    WT_Rx<=WT_Rx+6-RightX+LeftX;
            end
            else WT_Rx<=WT_Rx;
        end
end

//YC1_Rx
always@(posedge clk ,posedge rst)
begin
    if(rst) YC1_Rx<=200;
    else begin
        if(timer) begin
            if(YC1_Rx>=LeftX+8)
                YC1_Rx<=YC1_Rx-8;
            else
                YC1_Rx<=RightX+(YC1_Rx-LeftX-8);
        end
        else YC1_Rx<=YC1_Rx;
    end
end


//YC2_Rx
always@(posedge clk ,posedge rst)
begin
    if(rst) YC2_Rx<=600;
    else begin
        if(timer) begin
            if(YC2_Rx>=LeftX+8)
                YC2_Rx<=YC2_Rx-8;
            else
                YC2_Rx<=RightX+(YC2_Rx-LeftX-8);
        end
        else YC2_Rx<=YC2_Rx;
    end
end

//RC1_Rx
always@(posedge clk ,posedge rst)
    begin
        if(rst) RC1_Rx<=230;
        else begin
            if(timer) begin
                if(RC1_Rx<=RightX-6)
                    RC1_Rx<=RC1_Rx+6;
                else
                    RC1_Rx<=RC1_Rx+6-RightX+LeftX;
            end
            else RC1_Rx<=RC1_Rx;
        end
end
//RC2_Rx
always@(posedge clk ,posedge rst)
    begin
        if(rst) RC2_Rx<=630;
        else begin
            if(timer) begin
                if(RC2_Rx<=RightX-6)
                    RC2_Rx<=RC2_Rx+6;
                else
                    RC2_Rx<=RC2_Rx+6-RightX+LeftX;
            end
            else RC2_Rx<=RC2_Rx;
        end
end

// End Of VGA


//begin of keyboard

reg nState, cState;
reg [21:0] kReg;
reg [7:0] kData;
reg [3:0] kCounter;
wire check;

assign check = kReg[1]^kReg[2]^kReg[3]^kReg[4]^kReg[5]^kReg[6]^kReg[7]^kReg[8]^kReg[9];

always@(posedge clk, posedge rst)
begin
	if(rst)  cState <= 0;
	else begin
		cState <= nState;
		nState <= PSCLK;
	end
end

always@(posedge clk, posedge rst)
begin
	if(rst) kCounter <= 0;
	else begin
		if({cState,nState} == 2'b10) begin
			if(kCounter == 10) kCounter <= 0;
			else kCounter <= kCounter + 1;
		end else kCounter <= kCounter;
	end
end

// kReg
always@(posedge clk, posedge rst)
begin
	if(rst) kReg <= 0;
	else begin
		case({cState,nState})
			2'b10: kReg <= {PSDATA, kReg[21:1]};
			default: kReg <= kReg;
		endcase
	end
end

// kData
always@(posedge clk, posedge rst)
begin
	if(rst) kData <= 0;
	else begin
		if(kCounter == 4'd0 && check == 1'b1) begin
			if(kReg[11:1] == 11'hXX) kData <= 8'd0;
			else kData <= kReg[19:12];
		end
		else kData <= kData;
	end
end


reg sig_f0;
always@(posedge clk, posedge rst)
begin
	if(rst) sig_f0<=0;
	else begin
		if(kData==8'hf0)sig_f0<=1;
		else if(sig_f0) begin
			case(kData)
				8'h75: up <= 1; // up
				8'h74: right <= 1; // left
				8'h6B: left <= 1; // right
				8'h72: down <= 1; // down
			endcase
			sig_f0<=0;
			end
		else begin 
			sig_f0<=0;
			up<=0;
			left<=0;
			right<=0;
			down<=0;
		end
	end
end


//end of keyboard
endmodule
